PK   �j7Y#
���$  �c    cirkitFile.json���֑�oE� �.М�:����Hb�dH�O�ף�IO�eG����5�)�X�nvϐSoEFbð������%y����n]6�mW��moV����r�ڶo��?5���j]�6�w�������=��t�%����zǔ.m{S�E�P'��iRu�M�ICNy(ھ/Mi�/^-��@bS��A�`J+f�*�҉�
��b��)��A�`�T� U0e&f�*�23HLY��
�F��X"R J��V��X�%"��\�%"��`�%"��d�%"��h�%"��l�7o�m��VW����U�]�~J��w�ɋ� !ڣ��]on�{$/郄h��w��O	b�H!?%�%"`�,?%X�)A,)��D�����B~JKD
�)A,)�e\,)�W,���v�%"��v�%"��v�%"��O�k'�����ҝ�ҝ�Wn�3�( ܉C���Eg��x�J��I*?�9�9L,)��0�D��������s�X"R��ab�H!?��%"�|�/���k�򳈗����B>�KD
y�KD
y����8z���X"���ux���5��@�	��NX����t'�t'�g� uEq�'�	�	)�OHb�H��+?!�	I,)�'$���+�b�\��.�wB~K�2�����B���B�Fs�Ȧ4����er��#,�����6vP:�ҙ�bcg�����.N���s��A�K�6v;(a��������t�l��]�����t�̰�˰����Δ96v96vP:�ҙ��Ʈ��JGX:~<9;,���fp���m/�������G`>~l?������x��4�|��G����,��x�8~`ǁ�#0�9X� ��u`��K1��+��0\`�B`�2��+�����O��{,��x���6��`��ǫu���,��x�8~��+�,`�c��ǂ����|��?������W���v?X>��z:p����G`>^	���`���k���,��x�%8~`���#0�?"�X>��Wp����G`>^���`�����C?�~��?�8�����ό&#� ��I.�����@��/l_�|��E��������|�|?�}����ރ��/X>�q� l�<ؾ`�������,���M8~`���#07� �l_�|���������ש����/X>�q;p����G`>n���`��gF�W�z��A���ҧ�����j���,���A��BI�}���N᳣�~��`�������,���8~`���#0�a��~�|��R����W��O �� v?X>�q�.p����G`>�7���`��ǭ����,���I6~)ؾ`��������,���18~`���G��͛�ͺ[�ʶ�yE}H���ħE��jJ�ָ��S�m>z�����mg?�G8s�qיÏ���~�5u���v�3��)�9��G���ǭ=禍4�y7zO�������p�xa��8w�0�F�ޛ;^����/�{���Nm�xa��^a6w�0�F��;^��Wu�=q	�o�z���'^a��^�4w�0�F/�8��]�6�N�ͫ��y'a�O*g�PeY�s���i���Go���o������uOMCIQe&N@�ܳ�O2���kL����>i��p�$qk�Ҥ(�"i�Mo�"�P�?��&���&)��b޸<���;!�Ҏ����y��'?��}�7�K#wۤq�O!�,��NCK�njg��IÅ�>d��a|�۔��j�]\�{����`.~c�$�2#�А"���c�@B���$d��a�@B��!�$d�nb�@B�,�$d�c�@B�}6�$d�*����+۰�M�R2�e�v�x���py���+�(%3\1J��=�B&X�+}� N�2�W*�1��+au�d��j &��7��q��(%3\R1�긅�q��.}��`u���8J��hAL�ٸ��q��.%��8��;XG)��7�	w%����B&Xw�����"!������LixmT��.+d��q��(%�� c��q��(%�9 ��	��V�QJ�6���6G)�n��{�|��k�aL�:�au��kbaL��*V�QJ��v�Ǡ��B�3����gX5��:`u��+�`L�:`u��+�`L�:`u|���`u�īP`7�a��6G)�j	���+8���U�eURa%VS/����J*��<^ W�U��TXMyܸ �
��+��Fߥ���h��
k������&����(*q=n����+����1\WVRa5�q��*0����j��F
pU`\5XI���	�1:�K��th��f��*�.%ۥ�H�x���R�%Z~�\'�:�K��th��y���80Zҡ�g�ub���ThI���0��Vǉ�В-��Љ��S��S����O��!#Gv�v���L��:��t\�
-����:�L��thy��Nlu|�
-���+��*�S�%��ˬ�/�:�L��thy�Nlu|�
-���Z>����2Zҡ�5�:���e*��C�k+ub���ThI��׈��VǗ�В-�uՉ��/S�%Z^���`��/S�%Z^{�[_�BK:���Z'�:�L��thy-�Nl��VTz\QǗ9_�t|�
-����|�������k�*��c@'�:�L��th�W�Nlu|�
-��r�����2Zҡ��:���e*��C�=8Tb�u|�
-��r/����2Zҡ�(:���e*��C˽]tb���ThI��{���Vi%��R2_�u|���e*��C�=�tb���ThI��{��VǗ�В-�p҉��/;A��V�B˽�tb���ThI��{j��6��2Z:E�x�9������ThI��{���VǗ�В-�jӉ��/S�%Z�9�[_�BK:��;O'�J]>��|�����˂�/S�%Z�e�[_�BK:�ܓQ'�:�L��th���Nlu|�
-��r�L�ئ:�L��th�קNlu|�
-��r�R����2Z�F;��g:��T9ӛv�ʙn�s�Q9�y{�ʙ^�3U�t���r��L�3��g����<7�@ɋ��s/}�+���s�V�+���s/0�+���s/�+���s/�+���,>��ʹ2�,>�.ȹ2�,>��Ź2�,>�^ùg]L�{{�\�T���^�7W���^^�Q��]�6�N�ͫ��y���O*g�PeY�s���q�ʣ�{�ʣG{�ʣ��uOMCIQe&N����O2���kL����q���x\\SΛ$b�&E�I�\hz[!�	�h�ʣ,&���&)��bڹ<ɣI�����3q'g���(K��M�Ҹ3m�FE!�,��NCK�njg'�LR�������L�۔7�j�-.�}������uw��VW����$��$H�ч���P� D !3XaH��B2�E����`�!D !3\:����pB2�K���ڸ���+�(%��r�a��n�o���_S�0��7�
8J��va�`5�`E�d���0L�:nau�d�W1L��7n��V�QJf!���V�QJf����V�QJf����V�QJfYc�au���8J��/�c�pWRp�R`u���8J���+`�`u���8J����`u���8J����`u���8J�a��`u���8J�/��p��q�au���8J��Ø`u���8J�dØ`u���8J� �n���x��q�/8�1��x��q�/p�1��n�no��x��q�/D�1��x��q�/|�1��x
��(%^hc���V��)�_43Z��Vݯm��
+���r� �
��+���r��
��+���r� �
��+��Fߥ�QoH4XI�5΃T�:���+���9�J\G=1 �`%VS�b�U�q�`%VS��a�U�q�`%VS�a�U�q�`%V~&X��8.Zҡ�g�ub�五l���"�E:�K��th�Ys���/Zҡ�g�ub���ThI����׉��S�%Z^à['�BK:��C'�:nL��thyM�Nlu�
-�������2Zҡ�5>:7t|�
-���Z%����2Zҡ�5W:�U�#�tKLǗY_fu|�
-���8����2Zҡ�|:���e*��C�kub���ThI���V��VǗ�В-�Չ��/S�%Z^�[_�BK:��fW��$_�BK:���X'�:�L��thy�Nlu|�
-���Zp��*=������/s:����2Zҡ��:���e*��C�=tb���ThI��{%��VǗ�В-�|Љ��/S�%Z�]�[_�BK:�܃C%�^Ǘ�В-�щ��/S�%Z[_�BK:���E'�:�L��th�G�Nl�V�)-%��e^Ǘy_�BK:��3H'�:�L��th���Nlu|�
-��r'����2Zҡ�^T:���e*��C�=�Tbt|�
-��ro0����2Zҡ�g:���e*��C˽�tb���ThI��{���VǗ�В-��Ӊ�R��6:�,������ThI��{��VǗ�В-�dԉ��/S�%Z�-�[_�BK:��#S%���/S�%Z���[_�BK:�ܳT'�:�L�����|s��N�3U�����r����w�CT�tޞ�r�W�L�3ݭg���G=S�L�*gz>��:P�b���K_��`��ܫU��`2��L��`r��kB��`����8�ʀj0&�Ͻ�r�&�Ͻr�&�Ͻqq�&�Ͻ�p�Y����8W4��d���͕�d��}��|W���j�*�y^��h���4TY���>>q����ឤ��ў�����u�S�PRT����8C�|�̧��ӧi�x\&�<�ԅ�&��XťIQ4E�8��VEf�1���(��C��I
j��v.O��_�*��L���Y&�<��gy��4�Lۤ�@QH*K.��В����	,�T0,�s��2���\m���qq�.oW�����-W�r�m����ŋ��9���̊]�z����܉'�}!N<�p�W�Iq��B�=�?�q?<)��uܙN�;Ax�gx��R4>���VH����@z����mKOz��7D\�z��de۽��g+պ=5qyY�ƿ�������f�&�$B������c��3�O�����_�T����U(�͖�
����� �
}) �����;��|���k' *�%�!Td9�8a.�`@ Wv>��������_F�8�p��8&��H��cnW�My��v�����7}���r�)oW���$P|˱�!�%��r�b	3��R�%�p�_H!�0�s�B
���SR�%�𜫐B,a��d�b	3<g+�K��9]!�X���-D�D�O@�$@�k����R@%@�k����R@%@!�k����R�0��x!��GX©4��q�%4�P|�f�|��1yE�^����\��їr ��_���/�r ��_���/S�r ��P^�f�PB�;���\��jH9���ԙ	� �uX;r�%��J{I)Vc!Zr�^;�]���4x��,��z�9 ��J�\���.�J��f�wp J�Lu�ܥ�(�0Օkp�c ��z@=�kpW] ǉ�P^�ܼp����#��>���,|� �8��&�TP��4�5��#�P��4�5�Y �P��4��Yxq5 J�\���n�f�)`�+��` �����d��w8�}1����g�Q�;�$~X>�r�������|����A��#0_�.������G`�8� �o�\��X>��y 8~�F������ϔ���8=H��|�3�o7N?,����Z�$~X>���	4ځ�		M�O��cw!p��!�6"�v"`BB�Ӻ�����Є��1:�hG&$4!?%��!ڕ�		M�Ox�c�v&`BB��U����	�p�X��'��_!�aE@��̫�!E{0!�	y	�26�ŀ		M��/�1D�0!�	y�:���)�*hc�.Ƣ]��Є�dC������c�v1`BB�R)t�.LHhB^慎!�ŀ		M�K��1D�0!�	yy:�h�&$4!/D?.��)`BB�Ft�>LHhBs�C�O�{��w����/��_h���>š}
��Єf��*����蒬��;�W�C��-`BB�htѶLHhB^���!ڶ�		M�K��1D�0!�	y�<8�m[���&�%���m��Єܮ C�m��[-�c��-`BBr�t��V��Vжţm�G�0!�	�=:�h�&$4!�A��S���&4��A11|�0��cB��-m[���&4o��,�D�0��e���yB�.&�]��Є��C������c�v1`BBrG%t�.LHhB���!|>|>����	h&$4!w�B��b���&�b��]��Є��C�m��[��c��m��Є�fC�O��[�c��)`Bz��ټ�ެ���l�Wԇ�/*J|ZD���$k��>�����9�?js8s��=��񣮭3Ǐ���?�:s�����񣮤3Ǐ:��?j�97�	(���;��
Hsp�ַ��,�gm��4ǯC�+ ������
�k�4�oҚ+ ����
H3q�����L��i�9M���7"�����8~=�\i&�߱�Q��]�6�N�ͫ��y�j�O*g�PeY�s���j�����I�8���{jJ�*3q�g��}��45]c�4���I���ԅ�&���x�&E�I�\hz[!�x����|��C��I
j��@.O�8WO�����3q���I���>˛ԥ�m�h($�%��ih��M�샟?i������~��8n��{����~��pq�b����o�/�oy��0�!�_D������o3l�[oJ�-���[oN�=� ��G�A�GXay���GXay���G8��x���f�Z.�|���N�Z|ȟ4!�LI��S��ᾼ�G�v��ݎ�s7��>~�!��[OzG�q�1�ᚑ��cB/$�LFx��iL��£|�jiLh��Nج�x����0��{���px	�ʟ�rR(��~��2��2)��%YΝ�ʥeH�z��u��j���qW^Uuwť}\��v�8�b:�ʎ��~�ǿ
w�
�_��_��һ_��_��_�񯲻_e�_�w��y:S]]����Z���ju���4)��+m���mWf&�8�+o~�]}�z�y�I>������ծ��n�����u�ݭ�a&��z�p��H�춫�w1������\�P]�������o��yj~o����*��"�����ۯ֟�X\���My�m���Y�W݇�m��ݮ�]�y���c�Z��U���vۇH�ov�/Ϟ;�}��8���v�Mʋ̘�h/mf/�-ϳ�Ol�2�~�u'zu�Ɖ\��8Lk���]��:t]�_�G���f� Z.�zW���ФI�r�ٮ�J��]�^��j�\uwG�E�e���j�"-�ɟg����=�����_��ݶ�͇�YЅ�p��v*۾�nV�=�w���-����F�5������=:�|쎏�0r�~S����_�e��>�(��_6W���&����<���w�|�9�7�$��?2��c����������-/O���[���7u�}�U��y�no�;����_�e:��Y����L�Z�����I��Ժ"��/Bfc���&uU���.KB�Bґ�Ϛ�	մ/��t�Eؗ���N���.¯�����!��9�EO�E�gǹ��JjOr�S{\���=��SS{�$����/`n�ٶ�]�7�y�7���ֆ���S�����5m�7I�]�]�%ym\B>kMm���LJ�IWݦ%M�u�x^��(����r;i�t�Z8T���r'�{�թ�>���7e��O�Nm5�t��*���'i�I�w4I�Lg��������f��9��8{Nn6ʞ�[����V��9��({Nm5Ξ�[����V��9��({Nn5Ξ������V��9�U��Eq�gKN�lE��k�K�)�S[���$�[�S<�����s�������w/����������ݮy�r�|�X��Oz�ēEm3\�wMH�U�Ic߄,�s�a����M<����՗����)sk��m��DEg�uҶ����\:��Ͽ7.��ml�&�I���8.�\궢���8��0�������`���Ln(�S�9M�%����V]g��*���w����7K�)����g�{����U{_ٸ�O=�وD��g"�	�k]J��M�A(>������n}O�c+Oy�8�E��6)<�Ia��R��oO�|~������}�8S���Ӹ.��4�ǵ�ϲ��:���~��SY>N����E���<��C_��^�w?��~�^���f}�?��&���f���m�������/�]����Dv]���2�]V��Nr�8Y�������b��t��k�L''�&6w>�RRu}��!��En�������&im���$�)�Ivt46Kc ����4Y�
�����"):�'YSſď����k�}��a�j��t�����g�^�\?{���=�����v��g����ݶ[>�m�mo��6q~v������1]m6�u�T��	�mw�U�����؞���kvC����2��������N]<Cѯ��_���J{�bQ���?��.��}gm�G�8�*�v�=�i��ĥ��Ӟ��?��>��ys0�� W��u�����5��<_\z�.�|mm(�S���H�.O��'8߻"1qj�c�4�u�WaR�Lz6�8U��~�)Ť�p1i.\υOl�X��͞���%`s���_İ:~e؇����?)���ݽ�?+����^w���r�|�a��|��ǣ�?h��:U�k��������~��{���u����y{8���/Xj8�ă��}�ZߝUEOw�������a�A{[���Q���N��g|��Y���כ�z�u�{=������������Pn���/���.�t?#y�婭Rs�ի�q*��0(/>{��	4����K��A�8?7�I	p�Uv��?0(�&�ѣJz	?ȡ���8<�Ŕ:�n/Om51TN�=�?�?� �S����l�'�T�h=h�� �ীS�3����s���>]������p�̈́c.�'8��N~㏷
�J��|S��{��W��:�C�,��~x���?�����ǩ�{�V��j��]���L��<N1yR��qOK�ëbg�E6)-�yN�jb�zW���a����)&=���)��lZZ��l51y�8�Uh�R@�)!W4'�c�Dp��g�3י�)��=�_��/�������T���+1n����޵�ַ���͛/w��������v�?]��}w�lW�wW���PK   �c7Y�/WYp � /   images/0f73fddc-80bd-46e2-8805-d6b40fad9a5d.png�{�[���7� �"��
H
����!� --R�R�%��������'�{ݬ����3�|bf6LIQ�KNVRya|�z\��� .���hF���=;Y-88ʎ��.s�W�CG)M�W�&�.���p...��6���vƬ����{��pp�pr�b��;��:P7Ƴ�r�E"����Hږ�Z�;_�w�L���of%�mZ1f
o&l�qe��{��p�2x)*�|�W,�<!d�"�	��-��7��RA�voe;�YG��h�v*�e�É�_
#`���z��7�D��ފ�y��.JH����B����~��fI�wF������7�7���]�=r'�s,�>������q�`z1��f��9�6���d�ޑ�@G��Ig�t� �}��Y�1�,X!p�$E%!���s��#O��Hĵ��%���$��cM-x��Jcl�W>���VxeAKK�9���N:p�FĊ㈹��,��&�C�1D1s�E���Z��yұ����駬xB�єq�����2�WM[e��xf=��a�1�#N�B>��P��7�(�jA��#��G�����b�q*����-��	��$�կϗ�����p�Ϲ�R�ፊ���_�`���|��L�O	��H�űdr��٭�c��I�a� :7S(����I�Ӈ�7)�\�La-<U 7�󴪟U"X�J�y��3�˃��`��]��W��M���&�0����ԀԒ+.�S�h�I�63���+�&��ƞ!��W\j�L���>��p�+96��u�U񾧈���i޵�>k���L)��:g�����=�ƨ���UP.p�ړ�k�}�ASl]{[*�՞������Ǔ�����zf��8��H5��4@%�ltX�k>�"_�"Z} �גs�PV�p�m�l�1����i��g��eA�A5,.�/G������Zu6��_��dL?Yҥ�u���� nCv3"��@��ʷ���&�"8j4V"A]�<^AJ�"���d�����W�ۙ�-�Vy����ș��M+>�X���wij���y����Q��m�(M￱��*R�(�Q��?~z�0�U����7_W�&��fW�gw����I�Qbz�Z)kX���F�r8��{~�X�}.�4�Ī8N�ٕ̒���۸�n�����S�"��q��>n�hQJ���(�]�<?O;��;��:�G�"HC�oEr�6>Uֿ~2n�4n�t\ZZ)[((>�p�=�1�.��h��|'��6�ݎ���#�u,�gT���X�� �,���0�Oo*��Y�dZ6f�S��!6���詔�R�r夲���s����e���C���'z!S�Zj�xX��b�H��&F!������4�g�G��%�������S�� JT�M�3�r7x��A�>TQb�Itr��Ug��w��G���e�yb��ý�*LI�w����Ќ"3`�^���;		a��jvW=��T&�g}b��Df�>��%�C88a��C�� �eΝ������ko�1�W�W�s�܌���w�2��m���=T�N���5�Cw�h7�1)%	J���#%��$��8p;�,����B>���avHXx���0$E��[���*]�p���4	�
�:;��i�6��P�n\�px8#-�FU��Qs���WT�$b��Ý\	Y��VH���>��� !���^Zw��y��������Wf��p�ؕ�!hA� �;o�����x/���\���^�$yA		A�%�U8��������~m�U.B��ၯd1ѷ~pWޕ�4�����s�����M�l��M��eQ&rq>riv���媦o~9� lKKG�(�J;�1��P �.�'{д�hc����2�ms~�Im�I�S+k��:��O�1yL���G[H��,���(V/c�D<�DYpam�8�+ܽ3^��� �������2����L��HZ�����{t�Q��#-H����	�s������R�-Dg'Q阝`Xf��!���V���.��y�>V'��i+���W��ԸS$����jj�,qýJ�#s~�R��+�^��5c�
xi&�Փ$B���|�`��n��+4�,_�9����xQ�xс8jD�yLfu�����Q�Uv���n�)�]�lώɑ��c�{�*��1�9H>�~��n���t��۠��)U�W,q��?w������Ls��T*��<m�n������@�D`oٴxل�O����AR��2����X���T�hl방�f,u�@�J	\�d?��Ƃ?�'Λ�rָ����K��-���~q�'R�,b�X�,�?��v�ׁ�H��0��h�|?uF����<���ۛ�m\[t�l\��Fe��	�Wퟩ�? w��:c��k���6��+%�ߢ���Jz�1!��~ܵf��Xӛ�@]�l�@J����R^R,�-*���;���ݽ@e*e%�n��fݬ����ӻ�����N۫��P��o.y���`#V9�Uq�~bo�� ?RH�ߔ�������z��0�P��`x��C��ҸH`D�^�g���ٵe�/�~e)�a� g*f�����b��UYUߓ��y���if�F���"FP�\<n�7w�����5��낟��g�P���zA�a!"K!�P������<	R��9_�u�c��5�/x�2]�q��6�;�ie�s�җ�=a����r�Ъ51G5�4y?U�hѕ)-Q�.Q�#V�=�;#�Ϲi��r�����S�(ų+��}�+EǤ������a(����)��8�p�kDH�������!�r�k������:w�-�!����R�]˾"K2�Ē�ľ��ڦ��*��qr���9�M<��|�˕k��$B��(|�B��9�j���/h�r�VL��v5���� ��5����O����	�q���v;N/7B&��U��D�T#��-�\b��� g������ݲY��3H��+&�ke�,W�*���8y�ٗ<�j�TH
T�|4ۊ]��~.P����0UHZ���{���@�`0(��\�A�ML�8�ܓ��6�v�J�嬉���e�wb�J冾�#���ɚ�f� .쐮�Å.vLU�����V-S������ᢇ��{�����V+}Y__

p&k}�;��_�j0p2�D����Q���zW��d ����K���F�)O�)G����-gb� du�}�xi?�ݿ�D�~t H� ��Oq'�UoO��>��z�}�A��ġa���w�����l/�n�[���� ��ߗ�f\�o��
㉒F��-��f?�e�BN�KM�F;*���F�R�Z΀P�E��T��
�?�~�8�A�@�P�x���[DZZ��tg/r[\�����/���x�2���a��ϗ�c�_?�h�V/CV�aB����0�[�Md�t������D	�g��V��q�	��aՀn'O߱f�DiS�	����b�m�H�~�p˲�qfH�1�[���Q(�x�c�Ls�f�u[BGD<3WLB)���h��_;�J7qTA�v��Q�O�ĩq����|+�������~��?8b9Q�DU�\]�l��q��ze��-�6! )�5���ˆp��"⹸@Z�O�� '�R�`�]	P�'����hY��/��J6�G7�(3�ԣ��;�"�SF$�盜����0>�W����k���J;��Ĝd��#�|x.h�H޿fUѲ&��q`���Ck[�y����Ռ}�\�4��["{Q9�����{������Ǣ$�	B:*�Oc=H�:^1U>;Ȗ��B��n�_~yCQW{�h�=mE�h�&�d���?*ʓ.Ś,!�ݶ{ར�U�=Pc�Q'�����0��g����� ��N/�YQ�^c���5��]%D ]����MB��g�7�q�`�܋���<w�F�q��G�F�H�1^@ka�rEc`�Py�lyҙ�e�[#Np��z�4�ˤ�D'KMCG�"\�l'�v`�߇4gS_P��[nmec%�`|�莵l{��\{;��x忉9�s�=�	���4�5���,;U���%Z�Z�!S�'AH�k�����uhu]]�{�����2^D7��`d\\�Pז� P�]�dc'���_Τۖ�JF$@�Q��[�uԤ�^���^ֱ��"rﲽ(�� �T|֭4~:����~$Ӭ~6iB���=V����u��^^�\&����{!]���+++������@˄q���XLO=�L�-(z!A�W�&y{s�������@�ܮ�|6��y���.�K/�P�ɶ��ڃiy��]n��a�j�2}kk���2M����H�SӇ,v���=��rj4����3��(ia���j�Ȩ(}WW�h���M���*50����OM����N�����5j�S�y��2_���<dD�v�hSۧΈ3�3�$Y�i�D����toX�����ATL���u����c�M�]�9���E�ӣ��&`��<�/�����	�*$�>y�Nߺ�Χٖ��"�桥��v�������u��000�|��vY��M��*�d2X[G��#��%�;_��p-���K�qr�zp�1���x:֤���@a��C�v(Sqt����Sss_9�����+p�b�4��SC�&�[�TI�OjM���3�J�<(w��JKNj�Ə�w�w{���JxQ�֯�ON^AA��]8{x��D)�N`�Q|9��S��>T|�ӭ�j�	��mE�	�
���?�6C�{x2	�>z�uM��Lv I�r%	i7�9�]C���/Ā�z~��MJJ����W/3vҢh�?���`>c#v���@$Nh�Ť�:�f,�$���yL�x<�X��-0������Bv.� :�h�q��E�3w�u^Z��>�Z�$��.����o��ώO�b�D��w�TK���Tֶ���.ʤvz���u�ϋ�mM�/ �҉҉��?�[�*`�T��!�1��������� }�JJ�?�s�v,}	WS�s�j�ϗ��S��z���D��ړ�ţ�G8����-W�
�I=�F��1��L
qJ�%2�Dv2ސ||�06��}��
9�!cܠPWf�,����o~4��8km��<+����������z�ۗ��ښZZ�p�"�	��gi�T��j�0G~��O������Ԙ ٬��I�z�jB�R�ʢ��>j��jh����P�_q�?�bJǚ���-����D Z��L�ұ��ki�{@K?�Vyy:_<HA�C����uF��lRl�b���ǰl��L���"�U���4��b�%\��qt�����-���ٯ��Q������a:�Y3b���*����~��]?�9����B��F89���7��VЂ$RR2|a�雴B��>C����#�T��֦��1;^��L��*ȶ?50�4�h�+�k�bR��Hp�����	K'��ѹ�VD��� -g]�*��፥��H3�� 9��0�ˣeAz�����3�b�����DsL=,҂��|�,��|�羶��sTI������2�| >��2����N���g
?gЛb��X/�<_��7�Y!M��c	B.���75�~�A��r���Y��&}0O��丘J�����Ԭ�l�kT�4��@�9���J�g��711a��I`|yre��� ����̙���Rk',�tm\��m׼hm�.�4d0IT�u|�����T�f���A���J�6uC�X�r����ϊaօN	���₟U�5r �-_���kx���6���u��W��_��~ֺ?-<dcӱ�6�������K�%�B�� �2����W{��"�r�v�_�2���_f��lny_�{?�&�.Ƞw�}�Ue�	��l_Op2�%���}�ٌX �2:ե9�.U�L0��JE�u�*������5�G��ɷ?�t���7�y�FO{9rU����dd�̄Rk%��3ADwŇ�*�0$�[X���@3%~x���c�e��I�=�N��dG���1BФzv�����놬i�J�Z�������I��a�'ul���A�߾��:48$�	�,�"o<�pW�辒��A=V�pMm�D��f�7N�*����ףA޸Ag��dR�X�S+ϡ�}���^��˙kU�?�%�������+x����k�&��^�T	��m`3��R�ΘE���%��.,֛��zS�����;����e��=�������I�p�I<�}��;:S���3._Ɲs��ӈK�Cy��X1�%�lz=ڶ-A����G�(JK�N���/(Oj�م��d鿏y�E��C���"�22<<?�������{��R���i<Ƹ�S�z M���� �i��1&&��.?�b���QT��}cSkv����\�V?s�	�2�s�W���ys��y/\<boW�]�?��W�(j��	�u�cYixw�T���F��f?Z�6�
��ؤ�R���M�%�ў�2��:ۛ]�@>}:Q��>k󦘰�c�����>X�%+1 F� x��ky���4�X�˕�^������mX5q8����FC;�=p���V47?�K�>�ۗ�B������7f_w�!��Y�B%0Õ�9�-û��x�>?^���[Z
L[�cuP��ϐ�_l+ ����$�8�፦B����z^�OHD�{�?Y3��v�qo�������#�`z9�	Ew�K�0�VN�>���w�T/��}-]��wگM|�s+��3y�p�_��{bh/������ O��u�4��)Є&榧�}0�X�y�/,�$��J��i�������5i�k
\δ���/�N��&\�U��/�ޙԆ%&>��i�j��~U���l�P1h�A��<郿e �+fG�Rz`�z�J�ǒ�;�g[[kC���ݱ�l[�]nPĩt�r����>z�@T��Ͼ��T��]��q�C�Zm����s�hke�4���`��_��d>��c����]4[�@�kr�ϟy�s�L᡽+�	8�Z�r��>�&��
SS<�*�L����լr�.vy�E�jbJ����_�=s���l�9&*ƩQOM�ÜN����;<?��11���Gu��;b��!���Y���X�N���ϻ�mX%�շ��O��Yu?�N�z��8C&G-�F,�r��/�4�
�xf�&���}�GI��X�>(�I��Ͱ��q'�cwP�u����e&���Y��$�o���C�L*�X�/�-}K�r�*)b�緘i��&��2�k��ѩ�uyp��ݢ6������/��<�����Л����%�#>�\�hE�]wF����Ct`�5N��� �l[����l(���Cv����\s���۬ta�pn�P�0��5��5� =� _6o#1��F:�C���"Dd w�&_�$�uy';�+�����%EY��\�M���L� ��-X��Mo3A�V{�H��O����l��َƦ�7�%b�5S�૗���������dZ���&FwŞ[S�JO���i[����X�s3P��������|�c$@׷����3�����R��Bȝ@Bb�+�!!�	أLĈA�K+��/e�	*q���Q-��Y@�w�e.�j"�"7��H\=�Ŋލ�ؕqd�+�7Dͣh�_���� $��ȯ�C�.6w?���ݾ�m�^���^�PU{%m�F�D;S�߻m*������6�Ěw,_����W���ڔ�G�xh����H*��߁�khhȠ�(,������?!�E�����g_�M��z]���G[�RLM��]F8�Q�w�;���� �}9���]5�M*%w��z<���cM,]�0�MB�|�����/�Wꁁ٢1�N&y�7��S[��[���ݴFZ<��LYn�$B���p��~5��0O\257�`�u��MZQ�v�Hƿr�ݗ�;_[x>:�������J�0��~�0 �Y^���a�c���z����́�:�����z�c]��@�Y9��|7��1!��:2�ɱ��q�˝Zןa�,�G�a�v�x:��%�UU�&��#.7��m�>���'t3�%	J����A��f�7e6�Xoa3?�{U��{���'��4/^�R�?Q�5jƍ��8A��k�{������������/� �Uj���}��<���z�Y����z��N/M�iNb�O8Q�=.��\��r�
k��jPOn�!��X9��P����*&��VE���ֱn{%�=$=Z��mhй\�f��,x�m��m\�c������ti�>�]���)>���� 0��3;��z�Fb

�j�J&�#Q�P�e�/�{D����F��� �igǔ��ӂ�k3�^V��J�vt"�H�nK� ��3)p�7��(w�e�4�yVS����r��&��\���t���/��/QCw����3D�H�Z.` wF��L��[�3N�� ��y�7Ѵ�I��̮�Ψl��2l��RA�,�R�~A���n�UJ�LTA���`��bߨM��5̇���(K("��W~h����ږe^�!�#n��
�eW��Δ��6|�a��J���oig�����m�f���"�@M���k4Xӻ4�h�6̉*��|n[����`���
��ɾS+������"Q�v�����-ЯO$����2����q�+|�����s��D��u�n2v�ӻ|�P~�K %�.����K��	��\��Ԅ��hQ�@�۠_�˅��/ޘ���ʥ�=i�������sB8��\�'�+ %�<��c�����N����O��2[�Ώ�@(%>W���B�6�wv��pW�3����j����Z��h�:��IGHˀ7i�[����֖��I=�MG�0ɼ��uXd���Wa�0�����qc�FS���,q���:�튠3�����::����wS�E��q����w'�ǼU���c��
cv��xB݊�i��{z��c�՝���O�p-)���?���󃆨{]�eӳ}�g9Y�}gE+t����o���))�Sj�RJK�7w5��>M[�d�I�����%���^����4��ƛc��2�˾a�9�9G�s�BY�mx|I�!��5w�����4�����s�lQ4Wɵ��gFЊ�p���ȤI	��.�v�1���d�n�y�k��~��$�(���m	���Xޙ�u�9��a�@[��� Zl
�N&&�ۏ���h/U�a�����h�p������q�;����^2�q��zRǈ"�SJ�2E1�G@��鴆��^̜�44��]϶u��:�tGg�\���6�s�|��~�V��}����Yם��������F�Iޅ?�WT��
Mo�����*r�7�~,�gsx��u����?'��x0,���x�/z���˪�F�R=O=��Е�:����s�������I멚�P�k����{�ffŖ![��Ězz�M����	rwjQ�R�
�lZ�tGu�_;姛gǴ��xRT-���>&z�1�p���ws>u�[����4�_�)7��m���/k\��L)��1���!��'f|�-�N��Z�L���ãٔN�ӧO����n/&�Y�lU��4I �\Imb�ЎO�.��Ӭ5eڌ!�zr�i3����Dud�)��
sRuuu��9EƳ���ҿ>�=����2�퀝���E���j��k@q�'�F�Ń������:^KK��ز-��U�WMt�^�<,��l�L3Eϗe������S��@j��ܫ���m���1���um��uS
t+��_Czrs����V�/�Mj�'�qZ���3���#��a��o��ٶ�3d(2��(`u,��3=x�D��u�Op�����N����|ʈ�"��Ӝ�+�Z��V7�>�qi��{98��5kg'��L�9a:��0��.��3�{�Q tUJ-���O���3��FY
T�����n;��ۣ(g���
�M�Q�܊� I�߆���)?�Ͽ"@���v�Ȁ�<� ���!��~0}`��e�Ϫܮ��H��5�
EA�ݞm�2Ĉ�5�~BhQ��ڱ�&��;H���o��ݽ��Gt7�׽��ߟ�JLeɽ"��%�Z��B�G{�u�s:�r#��w~����m�4�YJL��v�s��QL���
���Lܴ�\�m�`��:N[��.,�����g�)�ˬ/����TW�7�c��2��E8{�c���9��e�$I<˒{���T��m%�|sG5�=�+>�pm�e'/H3EW_�½�3vz��"��v{���ا�	�O�rY0�����Ɛw�}����_�]n�V�]5�]=��:l��¢��Gl*d(݌r��=�(�g;����P��EUgNdYLh�s$M�r������P4ˣ���߷��#2*&ջH5��J��L�?������������1睊D���t���iևR�����f���jq��Y�k�9����E��v��[-���(rn���}����M&�
)Qݯ����|��K���N�]Ȓ#?j�G#����'6��2�E�eO
i��˓&�_��4LDKK�3 �����yL�q���7o�e�y��LLE�3���j$�IV��K�y�D��|Awѿ9|b�jbA^������ˀ�$|���۶����x�}��B�K��'���K�Iu���<���zzzZ����A;��D 1�8a,�5'V��G^M�I�|,XV�צ���S��{b��r߳��@o!�f�K��%�t��ɼ�>k'�����p֊�9�{!�qE��j�u�Q���o]8��OAu�y�5Jp.����J<�m�(������]I5{;˹��@,e�lCo�Wm0�=����^f��3����9 �� b�k|�t�;���a4���M�z���xf��C1�]�����X��& ��5�.���r3G��u��Ϗ�v��98�/)\�����ѐ�fw˷�.��o�Z2	�4bf�z��?GE�3�G���rV5Q0B�G�2�	:�A����di�N�v��X��≝_��J≔2��e:Y:�1F�o�^� L\�ʲ$F�c�N(� �x�'BFF&�>!^Zڹrоr�	� ��=Yyڽ�29jœ˄��, y���b��վ��0�)����<1�AQ�B�0�nS�共���s�p�j����ul�*D���(��\:OFߖ������Ml�%�ܟn�����pᢡ�CD��~f�r�a{�+�ٷWи>���+�� ���=.4���{1����X��!]�r�o�Q!�M_��I��qX��T��4_�&m�s����n�~v�-s�I��V�ؽ��y���'%&��+< �F̀B�#���P{����
�ta���>�����Ĕ�^FC��������*����}�/M��ن�N�^#�U��`%�����¼�M���|B�FD�����,?~#q�������D��73����_]���ZZl����-P(s�������c�����3�����Ń5{�7����ߙe6�M͍f��k�'��xH�g�7���ƍG��#ߪ�1'�3'�4E���ض];�9�/FQ���zˣ�L�vz�l%f%!��h�-�96y�P���VS�8��z%|#��L���zz���S>D��$ (�GM^?�ߞ�&�`̒�`	�L5%1������O��ܤ�����_�媗�n6����q=к��)[����%-Hyw`�k��VӤv��z?*5���t~�� ��XN)s�2h�9���7c[�{�q����p��m�/�Xsv��eh�0qp���ŕ	�¿������������8�..vH��7��ʕ���&&���D�:�|���0| ����=ŗc�]��m$�	���M�|��P�MT��"��$o��2|`�_��I������X^d�����x_>��O�`�oB���AZ�Z���:ME.��>�9���D"���ܳ�V`�����]H�m�v�HH@����9��[�Mr�ie��]k�ǃ{@ ����F�S � @��e��3 ��r+C�+�?�1��B��d��n���sd��2fe��@��]�<J �_f���>ӻ��33���F��e�ϻ��ss�QKgv���;nL2�:ƾ��JX��u!�8?z�לB.�kL�`�[��O��R�<�I��8�%�v��嶻�Lv���k����y]�s@�r�׈���v�)m��Tg��.O�������������Z�\6qa([���W��qtt�u�U3��g:�\l�����5�����%�Q��C<I��E�~��&c�FSHp����_g�lG�x�� �[�D8@�:Lj�==?[:?�c��X��~j��>P�*/t׎�p��3L�w$�m{���!��r���T�Z��;�h���{U�2�?:W�y�`�x�i��������\��G�8jj����&��Ϋ�a2��*`>}O/�򥡑��m��69��zѩ���/������kp?�ЋV�����0�����K���R�k>(p-��ZY�E���
��F�-�vN�I�1Չa
�!ϲL��N󉾽}��K!q��'+���<�}4��c�8��b�[��G�V'��4����.��!.o��s��ھ����Z���,���0V<q<�izz����u-Q������FS��d�2xq~��n`>�Iv"�n2�o ����ڸ���'����:�6���c��׋��՚�`�<^���N��4�P-�h�Le
�7��;����EQVV&4{$v�߷�O�J��M=��A��5,�M�k��jE������G�����X���x\�1�qfHϤ$6㊖^k���p[o�y�4pY�d7�޵�"\�Z����V	����_�y�� ���C�G�i����َ�H�Os��4\��wtttH3����ugݙ?��i�1�*���x�j�ѭ�j ޹�n���������y��DYz�_�YW�{F�Ӹ�Je��çm�`�uXQcz�i���^_�1�S����v����f�N�6��X�i�:�!���IIIwf�,Y`7:��U�	dq8N����l7yF��3��o�.~8�Bs��R𫩳�[L�L�Y�aSJ�>�Y֑��y�L<����ʜ��8�]�z����Ra�:�V����[h�?~�������[�m1���&��.��&�Z=r�[y��x]NHHDT��8�r�O��I�	6�B���z:�_�TA�< �dh�©j�L�ٹ��m�}||���D��Pi��?�lN[��E�~��)-5�3�T�ēy���>#����Գ�?�/$�oUW�\����1���D�^��-ߐ��V���v[�ɦ���o��)cxD�Z[~�AB�E��q��9�M���^�t�u�KPM�na��2����&7���f���tc���L&@G.h(��U[O��T0�LmŜ�ˌ#*R̬�����-��/��.>����gX<��f&���ӓiY�w`������w0[Xq��{jj�WG 11�>��a7s�4�wP��w.ۥ|Z�E]C}������RA��VN�$���F�sc�O���d��L�/]���ۛ^�덣�?ʯ��]�9��ύn���՗�c�
cU�^x��=L`b?���h�t���J+��u6���� p`����Sm����*yyV�ۨ��������n������^L����[*W�"�[��� O@��	��$ٹ���۠�fRʱ�&q���O�^Ը�+��՚����6�cD��D~�[�.�-M�q�ӌ����K�s+Zor�մ��&l�2�����s��6����H�U�6pb�E���
�ƙ��!��+ez�[Y2i��N�yhjj@\
-�97�]�F�B&pn�:��I̷wE�px0���p����E��!H)��q�9��������P�l�U/""��ʊ���	�s��������VR{PZ�7mu�2���sl�2`}�L��w�]����TW�K)�x�mn�Ԋ\�B��p��)R;�n��[&��?w���s�Ӟ5�cm]���w'r/��vMI�,��^���?�[M��ܨ�l5$}�����q�����̞]�f6S9��Ɨ��SmH���,���3]��
@�m ��$����:v����+����r;�XA�/�d�����Q��;����:�69(���CK-w3�D�I�K[�A�n��ƙ1"���g�%O c�f��N&�gt3�8��6v���N�I��
W�9f��St����~�*��؉�llO�%�9cH�n�����(��o7�L��b�2�x�Ϧ��8��a�(���F�:SR�Jz�܉Z�\���c(>��T`'�+��;f6`�Hg�p�T���g��#�D����0'����^�Ś*��;#���h{�)�{;BS�e�r��r��{�N���m�͙�p*��}f�*�8�ښ0o#ӢKu�}�cߨ����5'Q�*([4�%�zK��!�p��"�Θ(@� �O���[W��������$(�	�&��ʻ��.�ɀI8�uY��A-nك�I
��>�-U]�n(��ś9з�:�	��	K(zIK��^S�2�
=��1~���O��D�=��m(�>�Y,��7�?{f�D�#I ȡl��]pH�w � ��G�Sܠ����2
�m@���F�-�-U?/��]�����1� ��Ý��^<ٞ�����ʝ���L��D�*����_(�ޕ����ʻ=�U��-o�g�c�/��g��S��*u�������]^kkweߞg��旝_ʌ��w�W|ߪ(RI�P��#��>�3e��~�ڃ�Hd?�E���h���u��&+
����уLLn|N����Lt�2)8<q$x���'N8�j�q�6ۘ�7o�Q߸�d���O!���8���.���/O�aC'�A��
�������Ҋ�����a�'�v՗^ٯZ,5��ZaG�{�ɞu@Ek&MB=�����կz`�d�%,�=rg�ܬ33~���=�@\q���[4���Nr������
�=�Bϰ�W�H`:��KE"׏(=v��94��̴Z�OML�A���� ��`_���^�ey�=`�c���j�;���a�ɂ�� �{�Gh�J�6���O��-**b|_;������2Oɋ��(����A8U�������eY��1<~/�y���Y 7M���ވ���7X%���Ѯ��6��<.��N)G炔�g����n#��K�_���Mn����_4�A��d����I�޲���'~?f�����gJ��<��+
����8Hb�	%���ٽ�+?#�i%#T�J
�W?��+ږ�:{RKQM�ǠO��ݽ|]As���'*�w��w���<�L։.hCҠ���3���Dk��|���| w9���|9�cozlo�mWA��̓���f�E�������]|Jiii�'b��o$����]���?S�X�ɚ��(�0$G~�Z5p婩$`\����5d�:k���\jɂ�����ب��W=B�P�>t�ܯ�)��+$���\�Z		���!m-�Ǝ��/���m�g�����z�W�U��4��'��f��GĘ^:m�Y���cU��333��n�*a��ܱ�b/^D|�W5b'���B�̜X��ckcc��LP�����!/���0�C[=���s#� �~�c���g����g��܉0=�<�[�4mmvAN���6�\߾���Yc-���=��Wg�����!��~�L�?O/�U���T?U��j�����%J����I;& 'y����"��D�M���r��ڛ��w�4�)<T��1�M���+a�M�,K̷܈�Ax�[ʭ$�"#�glϛ��8���t.|
�>�%�����W#���/Z�d��=�Q�NP��Ζ���҈Rf�=�X�c���
�ZF<�T�RTKFF�R�K	�96���k�~B_ �*3r�΄��[rFƎ��F>z��U�`��u���Ƭ������X������H����~�Ѵ������X�	�<`֡z�����9��I	a�E�*T^&&(��>"�7�&#����DO�e��єP���H)((��B��A���������œ.ř*���;j�����𐓇�������m<oϻ��%���m0��+x��sZ�V�-��#T(�����j2U� J��� }��v�8��ˑ���=J�g۠�'�v
�$����0f��m��jԑf!��Ӊ�����U2��V+;9q|8�MKz�z����<u�,50.ݵ�B���N=X�VW�/./�}�	ё��˝!z��e (����k���Y@��&�QK�J��>�) 4�ƿ��e��X��r^h~ck/�x�Ή�UUo��5����^�.�PU�7>*1� ȿ�-�&�px:�ǅ�Y�^~��Ǐf�՚�I����5qѐ�aT�_M�װ���O<4䤘��`y�r��%B��rX�)���s�*��H6�0��szK�'�'v7����7����~f��Q���L�}y�:6�����Z�Q>a"�J�eOz����P��3��#k�3kH|���E�&+��b+�pr����ن��[a8�˨�k�?�����x��~�퓋�ˑn��"�1�IW���(=�Ŭ���(^�gzCj�r���7qO�	�zʍY�+�=%���*����|����d��k���&���.�H ����L��/.R��]!��<��A>�_��~Ql7��'�)<���d�����^�_�H^���|���T��n�ZH�v6Y�K���=�9��fJ%��˖|��YW��F�Uvf�iM��������a�����^�{Mf�ά�w^�Q�X�jlg�%�|�Y�԰��y$�7ʤê�v��~V�s��uw�Ϳ�(��t�1�[{����w�(c����Sx�
U7�"�m�G=��q�����	P�󿿶��t\�U�/��L` 	�C�=nP�yM��@�L�h�@w�(�ә�D�r�kˎ7^����.��3��������_�5�ۺÌ���SW�v+8lha��*�Kn�zH�W�I!u7Z-��(�,��_�蘭����ܱpʠ���w|��O��a*%��Q���ѐjxq��͎��!���/�Ul�s��"988���M[%=V�5�FҰl�ٜ�E7F��ו'�l����?�Q�PV�����}M����*��l�>%� - ������ ��)  - ]��ҮKwwwH����<�9(�2q�/f��õ���q�"���V�>��lO|�c�w��[D+v�g�Ź�"1��][)�e0�QXiẙ��s�!r�/{b���*�g�.z�G� �b�d�}j��[v�{'���;��8c�i)l	t)a $,�/i��4�}%����l�
�
VM{���k�^���׮��6gq܀�:�]��������ը@��)C?X�`���Qh-���L��A�S�W�=��e��CA�!a��w8fM�<i�m3ꜙh��fޅ8yٜ����{�6ϊ���f7��S,ߗ�u���ߪ�:�qJd�ÿ�V�/Ǥ��c���p$�A���3�]h1����CCC����qb��u�x%������&�Vo�SP
l���D� �7a�+��7�M9�/��.J��ǎ�6��8j�Hr���!��`3��WC��1�b!F	uu��q`\[H5 ��5��G�ϧF����QA���6�j�iP��3b��RP�2@\�D����.~��䞼Y7�1���eU;�D5��u
���T�e�����K��1�����&W����D����x+�:��vJK�� 0����X�WWS���CHZ���#�'b��R.��%��T'0<�#����:i;��{��A���qGې���d�ø�VϠrԕ�9�!��?��Z�K,��q3�j޹���C��vK�:��o��d��0�h��.Ƶ��[�L�g�E��| �iV��^Ìӏ35�3�Bǉ !�_U�ন��QQ�����ؽ�#gR��yZ�bO���&H��e�nWp��$�^D�q���[�5nu�y�_�� �M-:�;>h�c�7���P�)��_��˾�'��!\w���o�Ϳ��|�wvv�W�o4����\��T���a���~��5t�5���L�lя���7U�M6%%O��R���#b``��L=0qp@!�z��<��dxX���Mz*��~�g'��A0��������Lyt��щ��@g�w�8?`%�����~,HQ����16;؝�,rA��S����E��� �C\�3m�v��r�J�1��ӱd��n�@#>S�ȼ�+g��&������=%��vL�LA*&��kNN$	�l���?*��ږ�ܨq��9B����S�Y2g�H��, ~r0O,��VF���z�Ic��|Z�>�Uw ҝ�p���Y&s1��@?�uQ-�"MY3����M��Ho�Pn���ZmW���S����K�q���ϒ���T_�'�H�П~Y��/G<A�ej =-�,6Wj|~�d�i`(���cD�N�6��9�f�X8��MϜ.ό���|�o а޼ڼ�.T-���9�0ssS�c�������1�m;q�z��4��h3�0Z񙽣xj,�r Ȝ]��{Wq��2�N[	6�'JL@���݋Wψ�Ld��&Y $�u����J���X���De��9���O�4U"�n�$xR��$h��q`u4w�KF�u�A#�9�[������3�섨
�!��tg�J�.�6Riz�B�;7���?��S}8&Ws���m��,GĔ2�1�G�@W�%7�Z{�3/�i� 6���n��nc�6@�ܟ?�}?�r��l�o>�����H2m(ܘ1ܴ���OM�"K�EB_ފ���T:g����I��� a६��
� ���՟�CwOҪ����[�7��w�-o���[��;VR��`����#J��Z��1�f���,ŷ�o<�+Թ��蹲u�2gX���=�"��\!�Y@|��K�ucl��TL���Z�O�n�/��p�PcI/A+�M4���A�_K&>�+ȃZ��6�!������33<eÖb��L>>>�.-6Um��eti]\D���#���O�>�,�����EN�t6���6tɡ�,��6��k%��\N0G�b� -���ӤjI������kv������n��匡�]7^nv� �)�u ���g�8��x�����[6�葲w���� G�9upx.Z�� z��*�)��������)��1�+���YaW9�o?0��j��ʐg ];i!������>����,lw`o��y�c��?N�R�f���u��������u�Ü!��?aQW'K�  �E��\N���=��
��d��?��"���)�TD5�$�����D �ASS3e�ݎ?""bt~�� & ������mu�uZ48/~�"�`�诙�j[q�&���!yy��K:8��sY�sv�)1oA�D�R�>[�Xo���՗�]	R-�4�{�|%��O�XWW�<�4<TKm	d�:��q���-+��6[!���B�Ӝ-��b��n_;̱��`�I�p�B�!���,3�.j��� �Vf���!�&��M���;�.UۡL��y\�cʘ&F��hж76��ş�z�l��X�,5g��p�m��L���(�|�u���%:�g]==vv8�c7�x���<If�aļNg׭�L�z2�:Z[__}�5b��'`� �6y�����0��0?A�&o�h2�(`r�ߦ�a��X�0���	��c���t@Ji�#��$��.���܆��-Ur�Uh҉��yE"]�͘�$�/gv&�/@�J���v��X߲e�t��}U�1b�7 L�e$��*�?2�[q��3���'�MI ��rnV"R�t-O
Y����W�4ŰS5�G@#pU|��(�^�]����E��D�f��2�&#�6��<��݅j�Z�:PV��&���ȃ����?~Y�ϟ��AN����j��Eٰ��J����ԩm)���r��?��)&A�ƎE��<<������[L0G�T=Dh5�=n�!r�Z����축y��o@�#(�1�1{����׹w1&]���Ǧsk),���Y}���������	H��Ə],��G�.��6�83��RA���q罃8YB��1��d6����l`rf
�e����[q�\�G��84��q,qqq������p�ׯOd��@�'�
�e#y�T��q�0�j%�����N�Njh�K5��M�H�%X�]l��iի���%K��7Q��X�+���6���P� �Z�-��H9+T	J&^�`��ԋ���m�����Y&ͧ&�u�	�/Jt�N:'�醈�(��;ׯ���zǃdq.z��W�U'�$͞C�_{f䂿LJC���ƈT5J�S�&�����	��YE�����������JD����D���m����_�ˆ,Ȯ��@Ω��]�q� n>ڣ��
	�~��pkN����&�@���&�B�xG�[mI��O0^��dB���0�%�Y�K�h��=���pia���̤M:;&O�q��p��>mjZځa]GbVa[��wtKB .

j;$�fM0���mpC�F[����x��k�Xm���(lut��a˕C���P�~m��2oDK���h�v��e8Q��H��*U$���=�.�U�s�o!_�?�ٙa�HH��1��#Q�KjBA�i�9\������	,p����e�V���|zz�8�"������p`B �"Κ.Λ��&�GM������U�
�������G`с�,�Ӿ"�!� ����<�pb$��������o���h�S��q�t�vL�d�1k��� *�/�j��K��o߿	����Ii4.��
|��c&؅�'�],�c���3\�8�O�%���3�]���m�b��Y(Ն�,��>X��$���.{qd~f��ʽ�M��Rj����R�.��x��:	z��ەZ�^���#� f��dtV��V�}O*iA�����2PRRk)�NҰg�Zݝ�k0�hSSS°�	k:9�7����Zb�DZ0�R��l��� ��������KA���-Vz�M87ƴ^H������Թ��'l��:����r0I6���(�vL7��Mk�e�c Ոq�� �_z~��[�ZɄ�U6�ίpQn��?�b� O�z=�i��6�\�=yJ/�7�ݷ��yS��۠ڥ��S/�a���j���~= ��� �6N~$�q��bI!M?��d��E�j<�f&4o?������� ��TT��Ѭch8����^@�P�����U4B���x	+4�i�E��^}'��dcC�-����l�ӷ�lggg�쬒+���d�篈�D۩]8��sQ� ��$����4���Y�ZS��u@v������~߇����ˋ��Z�P�~&uZn��M 	�u4`4B\ L�����vM)�2�|z
�/+�3/P��+�M�Hu��
�H�����UԿ�
V	x�}L�fS�r1�*X3Pn�X����kǂp��@A�R�(�Yԫ�9����V�^]��_�����(��kc����q��������k��g��Y�ﶴ��?��*��"K������EP�$-B�\{��I]���7��	��6��e^�&"������4{���jyw-�b6�����+�7Yyv�#��G�cڋ�Q��_��F�#��Q��%�*n�f��u�c^Q&�p�7�[����:0�Ջ�i�LKK+�`gg��?4��&"�Kn��"��<�%R��Y�3&2��؊���4ɭL�[�����9��X�Ncvu�$Y/@0���}u�)E�f�[�� u�Y�e�R�t����9~�ܝ'"cv����\z>,6����V����[OU����YP{B������q��׃��Xo��z���uf�)��ȰV������|N����_�`��A搋ŀ�������5�l�m�z�v0��np�zF@��8ɴ�{�U�b���m��/���]t�������1'؄qG��P�8����E�0YY�J��.dkktq{��`�cU�l;+�v�-�O�e'��"����#Mdc䕍���B��� �!�V�$���%)��Z�O�%(�8b�b���c���\��ɩ�3��<�~mhMi���@�[��?��[Z�p^��P�au%b\�M~3��+ݙ�Ī��T!� `��ӆ4�Vu����:��_G�J�{O�9�1Ԫψ����RU|ŵ���P=cej�גK�i2�k��m9�B�1�ݗ�v�������b�e�<���*��$�-�4R��sX���tâ�+O�L�����bs100���)�F�
��V:��:��R�ʚג����߿�Qb�M^lO��j�}(������Y_#f(&&�����um�[��,%rnyR�����y�E�Ib���X���m�#5��Z�i��e�78�7�|�t2�M7��W��
D����8Y6����K�ie�X8�Y.K��7E/U�mlY���T^�����֕�5����4ӏ�t1�Ƚ֔ӏ[.ݖu�]n��ڹ-�h����ɕ⣊{ܥo�����ٽ!s9L �M�h�T�8���d���,$�$�Ҫ�;��z�MůZ�n��J�i~�.�D���YFz��_��& �0�5Lq�qn�3���꺿O�'�Tf$�l��O%uc<�F���x?����3�U(�(��\�*|d|��������B��k�p8��ZLYL�V�� /l�@b7�+�勢�QJa��^��`�?�|��'Ӌ�_��^�&��8CX�[{���Ie����:�|9�k��$��a�6�Q3U�<����7+��g���:�W���(���B������h��7W�3�{n��� ?VV��������%���XR�V��[��зF������3 ��I6�F�9K_�4Vsd3��lK��=������	I���*���n��a.��K|w�|�B���`��QR���H���M�RV*M-�0B%ef�-�U� �,E�H�� �ެ���9��	�{n��=�3�%G��a��v�'-}zZZZS27��4�C����6 ��#�kaɎ������3/>�5Y�����VVA�C�F�xh(�dcl�����Di4>y�I��	1��ӑWR��MA��(!��
/{���f�Z,���t�NHR,I�O�9��>ضe���X�����P1���+Ӫ$/�z6H�vt���d�`8�˙���C�/TB��G�T��Pa��7�Ѣk�ː��G�>S��~Y�E������C��Da@W�+)y��Ȯ=ݟH	�T{��8j��:���m)\�2t.�~����(�o:ɽ/�)�O�pw�z����:\��9(cǧ�T���<q���}�xOr}��챑�"�.pB�G��Cy�ڟd��t��җ��(�!��J ���H��J��9D��� <��E�
 ��Q�S��~�������W���^<��6]���'�=urB&++K�j��k��͢k�6�䚚ޅā���0���k�`S���#�y�f��}[��V��5���ֶ[�#�SbVg�"��M&�^Ҫ.*X�6��|c� �CּI1���9s�Z)�i����]o�4?�]M\�t�{�C����<X��{d����3����k6���W>�Hu������hv��9�O���ɇ�7*o�ɦ�x�A�*aIt�.�_J�u�,6go(}�?��%�c�{(k�8#�6�����O�r�˫��1ǣI�5�i��3C!��2�g��.i0s�T��?�nƵ��pY�
F�c�
6v�'*�������ۦ��U��LmSL��T�'_^����ZMJ
azz��_���6�?D��C��=����[��W�U���0~�F囹�]����R�[�o����y���҈Ty?g�#I,�+�g����^�?�zv�9Wz�z�s<�)���$ԱO+d�۠��?�~���:�y0�H�q7'y�g�KW����\��{7n��J�Ƶ3�3�#�^mp�?��jVy��h���1je�IN�,�j(��7�É��3���|�6LH��;<��ަ�N]��c�&��Z={��9.N6�I�����_/i(���%��;4:�)���@����2�����!�z��o	�|�0c�m���[��:�e�i��q�:��z�t�!�ӥ̾��j%���p��E���2�$���� F���<[`�mO�,�\M������_�l���z i��i3�&mjeʝm5Z�5y�&L��Oݐ3,s�.�����O���=���!�?D)�nb�8�Q�,[LM�G�����Qw�_���U�������k��?X' �gK�É�w��^3���x�?JQA/"C	�-�5�G�{�0�i�з�z[�����T;��2W�h����(x���L9���C���e��5T������/���(����}h�Ų�S���Lp�������/����W^�������� �9��!ݹ��IQ��;�,����G�G�6��x�=�f��R.�VH�?2�D����G�Noѯx�R�@!�O#V��WF�kB��՝K�Bm����βbl������aŦ���� ��-22��M�.c� �B\��:X�ٯ��;N�,A�囌~9i\\��W��z�	/]��-�D�2�j�º��2p- ��P��%S�{�L�ԏ�j3]�u��.`��Tۦ�˨�w�裭(ٮ�����3���������%�#pxJT��>ۍ�_0���sQ���#OA�Y�l�H�k�C�~�]�\�]�18�яR����^�o7*�����Y��>�?�X�뛨X��$�����
�+͞>���I�,�0�w=��Fuy����J�[�y_�H�����C��L��2w�����I�jq'�����O?�
Gۥ�C�cS�A'q�w7����j�������̅$Z��C���j7���7v5>�0
Y:�|�*�� ���
7{���w��䧊���)v�H�Wװ��:X�JX�`�O��g���0#���ŕa�756�����\z�^��-�co��×��� b9�)Sh�
1�ӝԳ�#T��O�alY+W
��Ӧ��z�:�5
�k�u����S;��>�>j(xY�Va�B������C�d��ԓլ�~��z{G��~�j���ɀ���G�p.�Ŭ�o3��sW*�(�>�L�/^�SV0��:NJ }嗺{�����~�����x2T�_�bKr���!}t��?�G�S�(����������r(o'�ɿco���I��z="����7À�$�����נ �=��'h<�g~���[#ծl��V(�����FQ�-�Wn�O�FX�'B]��/ sv%?�O�d�����9�*?� PW-F�^�C�-<���^����o��տg�2�����{pa�-!.�I�6��N��7��3�5�N�0�U\�oZ~n�7�:����v����\/R?*�6�gx��Z�6�.�k�kty%0�#�~���G3�n�`p-/���&Ҝ5]��
\Y�P$�]�����l���=?�BG�����V�B���ICk� M}��_�+C�0z�LOC]H��G:۱f�Fzշ;R���l=���?�k��4�����è_����Z�>�u>�s�y�K�Z���G�O��2��Ώ4��jt_���T�����HN͋ H�z�`��	�ɭ�aI��ea|\��vb����H�}ꄀ	�49č���Q�J�)Ks(D���Zht`I�98 =�h��M霝���k���J�F�P\C�ÄI�)����\�13iC�Jz��)��u�zY�m��$�f[J��wl��n�.ރ�B�D��W^^��{2�
޷�D)���#�Eƌ���)=�����Z��1�a�
r��aI�*�������є#�	 �%�ȡ���#HI��e�d�0 �Sm�1��K�#Ӱ��?t+,�\�������+����v�?��]��D��m��nR�{���#f\d��F�-��"��w��]�Bt��fy�?HaN�]-��<�F1X�Q�V��3O��q�� CS~��<e������q؍�
�N��m�9��^v�ά���ʲ�����@}i_�݌ӏ^��BA�w;U*J��EW�F{��N}}�ύ3�Y��RA��~4d�����T��D3�<�&�.-#�3��t�>����RdY���s�4#S���݉�����2�>dxX~"�E.��*0�
Vr(��bI�<�Ƴ���������*o2���&&�/g��X�bq�S7�����EQ����
p0�����#n�`A[O����Y�V��E�����������)�Z���|�p{�
�*<V������j��jb�z^x������������⯌�[�}����*���[�ԝx�eu`�O���Ӳ_FF&`ا��!u�:����]�K�Q��Fi���-���x���{���|�f� ���/Q�;�2��C�	���T����4��\����u�=:���p�b=|�G����z��@�>#�����O�r�3������i�hޗ�!�pQ�+�*��ji��`��.T�SmY��3B62����5g����c��G�W���	����;��a�Y�"���\��)��-꧸D������ �-��֡';��̽s����Q�O!��w$��~j ]c��J�3�젊�V��h{j�ĭ݇��F��%0��?�f��oUݢj@�z���ղ��w-R�1�ndϥe�^nњ=����|���Jvbm�: }�� f����tӉ�čzǂwta!&�����>1�r����	xk芑o���e�K�Ö5�� 3�l��:�=5!�uC�QR%S��)(-}��wtTy�aF��}r`��5���7�^f �{�q�>gggP,��jk�?���,�ri!HMK�gղ���h���:+ ~�N��$��l�}�x>{��p%��5M�QN^7�,��N��&�H�5܅��=Gцu�A���P���5�8�̥���e�NJ/rj��i9�ŗ@z��J�F9i�����M]�7���8?���+((4���@��y}��Tˤ[�u{�=E�+��$��/�asI:�1�BCC!������:� uΊY�E�1���||����]����4��+(Ky��j���V��Ή�b^�T�S*�HBK+��j6V�Ckk���,K�>��`�܇@���#����'�o�ު�<E8mC�'b��9�sF�QB�J=Y�Ӿ|�q0P���������/��=��b�OGq��i�N�a{hm��^�\"�D�k�G'>ЈP�k͵���/BND��ʽD��ֶ6v��ߺ�c�Xrrrє,888�1�X�Ϣ�>�c++F7�|M�@zD�w��fu�d�1����wX�6�0�<�#�	1����5�dtl,X,��|SH��Ê����G��H�w��!O��-3��f��-��O���=�ԝ�U,����s�`��݈R=���������fG�����&+�fw�(�6ʸn��%�2R|u�U�x7�JC(U��)r�΅ϭ�n�`-��%���"��������l��2�M?:ˤ~8�1Z�J3��2 ����&r/�iM�|z:Փ�@3FF�0��ݖmpc%�����e�=�d,/n�}��Z�.ϛ5pyY_&�zx�����݃+��� �ӡ��n���ڔ�x���?aLLLt732<<|�aa��H\
2
��⯺lMM����7+S#2���C���b���;_s�7��Y����Dw�Jwt$n����<�� ��eL��)��/;��l�y[��}����th��`�f�:����
�����n�v�+ɂ�4K�A�&�7'��ilܺ[Y����+���p#{���(��I�ڹ��+�Y*��8챗8�?�&�@<.��0T>i�8�(�d���զ&�0�UMl�Z�~S
`>�c����p�ʼ��w�m���eַ�,��&��U��`/--q��7�VB������}�2@����;9)�(��l���.=v�a�$s�N��)+���v�O���>̎3R|�mvvqQ�~����� 	�z�ᑑ�*,5 H�������j�5� ��:7-�/;�]�3R��>6����\��_�-!�1n]>9�n��z�ˑ.�� E�]"xE��J8Bl7dH��λ3ݨiױé���]K	��PS��� T�Și|:�MI�.H��3&xο[*S����ܶ*_��\Pe��;0��6֪e}�NfŇ�������������'�^+��RF��W�`=��K�ٴ��qp|h���(,�|��duX�d�k�*�j .*��_��U�����*�` L]L�q���a%%%��ūPc1��D56r�{�ª�������}�|�߿���N�[[^F���Љ�ňU^y9R��?'���7=##Y��_)?Q�)蚐�fr2�^�~��{{-VrlaA�)̆�P���E?�=�R�V ��ssR+Q���-T���{X��r�j��A��՞3�8�ا�u��|�d���E�a���i�D���ѫ�',�N_}�2�HRVdS��'NMVC��7)qbӖ��������H���U��a+����4.RxmB����]Ed�=Mt�L�1��Y�=,���T�XZC�2����OY���eڬ�Ŋ[�.�\�C���e�w֮|,l#�93Y�����kD TJ����4��0�+��m�M��R@&���_�� �X��D��P-����}��-���7�[��LME@@L��j�^�t�܋A	�%@�:ʧ��zyb���s(�t�m�eʖ�:������L	䠼�"Q����OgNNNH%:֛<mzMw�M+����^Ѕ�@x��3?�g[ӓ~��h��9������]�:n�7SE*a���Wb-as@|v�O����#���E������Z�Ӻ0�O���'���m��r>R`���v���	i�B��ߍ��Qc�fn��pQhג��{{%9�������X7G��&�6~}�QQ]=�[�/[�y~IMt�J<��sxW�1Қ=p��}��E�|�������{m �i�ݾGa�0T@W �-�;[�,A�C�7Ks��J�bIk�,� y��W?��mfD&0� n �y�X�I;�ߑ�>S������������F�,���K���˽	�A!��?r\IcvyY��(P��/s�ǚ]��&�*[��P�6t��>��x|������޻&l�E���k7Q��)􁆈CM�G`>��M:�u&�lW��ଁ�a����G���I��a�OȰ��F�6{b�e���M.P?<�n������hWu2	�>��.)N��������9
w��2��.��E�)�������666 ��i�a��m[3N#�x���0�4Ty�f�(3^��[G���у��=748h~p�:m�25I�0@���^Ӛ�:�c��JJ�6I��"���q�.��/E��x����D�(S��9L�6T�
�B`�[wx'�)o�MF[;\�T,	�n�ZP�)��ۘ��z�����q��M��	D��v@����Vw���@�� L��<=�МUԔM8`��T,�_P�Y�$�ƎS�l%U�ΘY���mB�*��!3�W&~��魭^���8Y�����'���KU���0�
�۰6G��ũ♁�*��g���:;v�k�-yI�v��u�"��HYB�C�f,���E��T>"��3����
�>�w=�"����BV�i�Ȯ�����a���1��ղ#~�,��Mk8XK���{���w|<pYω�7��
�-�jXޯ��.+�w��xw�)��w�hӻ��%�))�&�
ˀ�4'k����-I��2eMDb޼d��:=���5�z�8�\3I�	�pJ�gp]� ב���~ǖ�bCx�^cks��m�V��M���h61�x����*a:�rc$��F��kQ}[<�"�pss˞t��`����ȭ��i;��{n?�W{�ϑ�����!����&t��k����4�<kB��]Ħ�vj����Y�_�������ݠ�-�Ҫ� ���+��qR/@�$C���efB�G��"[�kx:V����~�C0��0�&(�U8q�.m�ۿ�ZMV��ݒ����ǻ�^)���h��W(�"5�pk�n�JH�*�XQ>+�~qM��Q�WU�&h�ҝ9u;:�>wm�Ew�B*W���}�|"�|t5��0/_x
%~�Zs򚱅	��j�!r�d Nj���2��qm˺����{̴6��W�?f�������x	ǝ�"�\�ZZ6�GI�J�ߐi
����ي۝��5����<%���p,�+������U��4��5��w]ۦ2>"2�]�S��۰"���F�A&���Al��wK�(7ď�� ��D���N��jo�B���V�M!��cZ��|W͖._�%��p�i�:�qĎ�<������QHw.%�e�kC�#�6�#܈�?��t��z����_2v�!��	E���㵅��b���
�:oB�T��1�uޑ�������c����2#���z����aŤ���mz$�]��q�}���\��*Ma��4b�G��Ҥk�GX���|s��\�к�~e�؊�p��4p�T}��j���G��C�� `ݥŦl��`L�����8��P����;�p �m�8`��͍�MEM���"�!�P\�rb�ʠ�ج���if�� P�1�n��s��w��������v����vmǉ&��{&�}�Q1j�N�^S'$3t�W�߾y���K�G�Wm}�9w\�g�EV4�w��d|:��X��Lq%���n0˧�J1���0��3�A��1���$H��;��`0u\&n����Okڮ�,��AG��u��6O%�ץ�v�F��H�a�����J��3s��Noǈq�sq`��o�3�I�Sq��O�TY��/2d�����)W �° �Lì�>(�2q;�%٢�X�Wx"h����(����w�]���ՑKU�+��[.-�(k?��m�&��=�Nt۔�ώ��S%x������u���9�5g�2N�p#�WOI���ֹ�x��׎կ�>Ҥi�C�m�~"~lK���#&Kjw<�tP�I'l\�^���`!�8����P�0P	z�a�{�F�F�fa�b�}t'�������O�d�G��`�#�*'Vtz�m{��y����7�֥~<��o�͛���V��gԪQ�����B��Q��Ӧʔ&�f�hw�P��_y���<'�:�ʅ� ����!ӻ���nM�4���7���.!L����8_"~6��pSt���YmL ��o��S��ż�љ��3ӚO[E�@�CT�a���H�-XZ��h*4�~`�p?�GW��u�x�b�R�E�������W�7�!�'<YY?�	O����OL%�<1)�&�{K$ن�!��Y�{�H�Lg
�Q�X��X����i�Mz�\�G�[�G�(��ѫ�����o�
�=�3��A	�"�Ǻ��\w'$$L�N��kܯ�	�6r�R��U×����6�f��\Nv
A�"[Dkx��9jt�P�ư� o�c�#��5���I*A̸�'���읳��1�Z\m�m���yǠ#�&Zֆ���\W�q�in�g��P�֏��#q��S�6�h&)9����D�����jh�1��8�)'Gz�]��z��}lY,Ԇ�~���[��%��ۏ}W�5f4X}:��Y���t��q��=��=���竕��A6ϼƶՠ�Sq���J��ރ��2��3Y��W��(�0�G9[���Q�D<Bh����f��J�&r�P(�}�ݣ�@�!�4���#�\�Ts�l̉\���m���ٲ`͑R-<;(s���"!���4(�4�2���T���	$B2V�8V&@��!����I�P&�*w������+��u�����m���.��Zy
9�&=�b�r�i��ؓwly����%9q͛(^�Z���jt��e<R�{~i���c�@��*��l�oa���-��*?�3� ��ɶ5�/�^:�,@��E��"�d{u����Lm6NaÚ�47i��%�Ѵ��-�}��|\�;��K	3������G�HȦ*�����͉�q�0�c����,���HO�R�h��[#��8�1o���|�+���X=�� ND*o̾g�Z������+R�rl�D\��-�!:���ת�,�Z�d�PP�����^���z��Ed���x�\��N��I!�e���w�mǖ���?��*ѽJ�{��7���݃�t�K}z�WVѢ��ȗ��R�!`�O=�?n���!W��"j�v)���%�~S�}�[@M��Pz������+�s�q	�V��zו��_{f��Y�Vw:�R|��o�u�W�d�&3���G�e�������ddc���o��g�-���\�ObRr(�ڿ�g�e&ո��՗�I��+�3�Ț�{L�%�zO�h��/��Mn�B�Cao��9�Z.��%��O+����� �DN�v"@�^��!7Q��l2��{c Ƌ�OM;t�/�XWP١p��a�A�DC����]ь9��!�2ޠs�جz�W�({h��w�y�c�W�6�SX�1����4���,ulu�E��ٶ�cP�a���|�N �k@W�>��J�����TS���s�k����
r��u�#'��"J�'Y��Ő�_����i�$F0nl��ff�&���l��.~F�����F�=e&c�C�_D�]e��X*���D�FQ#q��㝌ab&�տ�nwr��U��!S�X��B��e�6n}��R?�1�R52�W��Fn^���}^������+$���<���}Q3��������ڥ4� 9[�98b/�a��r �/��k#�0�"$����͊2)Q��<]��Ä��)�Ff����r�Z��b������ݞ$�:��6������`�Yv[�f,�+��H�`I�Hky!�	p��]�I�!$�vn��>|�x��<�G�ZajhW-M>4xR�d
w\h�))�,0@��+F�:��Ϟ�Tr�8����٣kw���l�}�#[�PEI�Sk���p	��r@@�J�EL|����Jd��w�|
��_>�@�[��9&u���� ���D|	��6i927��q�m͔�A`�Cz�$$y|�pw+D+D:��`�-��te�f�a�Q����E�:���V��Ż�į�,�hIV�u�,;��Xj�>�T��y�5��a�^j�{�D�A��U���I�"  ���Ȃr��<G�t��h~�,��I��e�^�:i<'6�y	�[�dM���G̓�*`.�p,YW�fZj�lLف�UbԽ�`����a]q+YwU���w�ڂЫ��"��>}cEz@똎�GRG//wHova`bJB1Q��I0���~�]�"�)Ր��PT��`��h$	"bdoa��7ir,$��X��==!����B�������R�S��k�>;.˦���Px	��Q��?PҮ�S�t���Z)�8��&'#L��qB�i"����JY�ˊ#+~Q\!�]�ױ1>��U3qq �m�@���\��א��-�Y�	*2N�,����bG��z��,�k�s�7�p�G����)�Ӊ��K���+d�FB�V�k)T?��~Z��_��g��O��3�%]*��f�<~6��A�7�s�ZPX��Ny����-�]V��at��ݪE|��m��M���xf���v�1��_���������<�,)��o�d��9�G��brT���ph<Y���u|��ۼS���N��k������x�2 9HNu����פ��~SW��~�����[����������Ǌ7��7��	�ZNL����*n��?��*TѠ�����(�)+���(6:V��D䐛'�
N|<�"L�m_3�W��E���vp�˗=���;�Mnho��Sepuu���W=�32���G"��,$���Y!v�{j,��&�B�FSda��>SH0Hʌ��R��0�:΃�i!r�H�Y=4��w.�w|k�/~�)�����gr����-;��*X}ӓ=~Y�W�{����5C>=�vu_I���;��5s���"�������l�D�zyE����<ll��B?V̀��'v��D����M&A��~�����)��9��X�C�5r��Z�� �����_W���$omm��t�!U��W @O�;�`��C��B,t6/���9�{��^�q^�UQ�a��))�&��Q�a��ǲ�lL���������%���������Ii�A@Z@:��钖�.��A��?�w��:k�L�w����~9�~��M���6���5ewg������Q+��#4�=��]wş)Q�eeѓI����gh+��m���ws��;oRg��&�aaS/�P��R�a��$�%ے��zzf�Ӟ/�� {-�����!��Ms� �a�h��.8�oa�6ĸ��爨�[^P�΢#���*�b��όq�)�ʈ�X����"�Fu�n�7��g�?�XD��k%֠7�7�@jϣ�8�n>�j\f�d+�ٿ�c���N��i;�:�~7ob�is�2{�!��;BBM�.���JL���]B��NP킯u������N���+ڼA�R�("

m���=�<�����;��RUƊe@q�����G��Z�.}�PWW��d��Hf���}(t���O��E��G<������M��*��&X���}����Ϧ���S������x�k4]��t�������'�"��i�hU�N]�gש�3tx ���9�4\"A�̕��5h!��gD3m_���}�-����|�F�w���8���$T�o7�-SC~���7�O��O�2*8[��j�X�Y8����'1m>�v����b�^xR���e�Px�Q�����;�i��gNn6I%�w&"!�oX�6�5��*llm�c�W� ��qt�;=�~h������j���Iy��2�%%b���|{ÀA�o �_F��2)�>Ʀ�377Mէ���Zk��ܹ���y��1�\ED�F��P���β��+�?�RZO �#8�����lP ^Fr���%==��G�e�y�I����bTa!���S��0q�;�8ߛ�ԉ��Nj�&�m��_&8��ɲ�]`2��24w�ޞa�
��m5.y�� i�vL�\��J����
���5g�F�r@D߃��&Q����%82�� �ɓ�w���_B�0�/%�pq*R�Fg����e�����^)����!�O�t�_He*E\^zx,XWT$'�w|�;�4l���f9)J��������������,�K{z�c��e��+"����6}�?�L�Xx/��T{��1۹�AG �(�s��B�:�0#VVV��(
��}''�3��l�2g�>���Z\aaa��Lk]�
��C1��Yoz7�n� l@�1�ޣ[p���ݛL5�y��D��]#J�lA��J��Jz�P�^�٪��N������(Rl5܃�WAP-X7mצ42�]V��|ѯF �iV�e����).�����K�p���ȴ��دp&&&��BA*4fᖦ=���"Rǚ���Q8���hQEo�B���g8�M�7�߿�L�<��o�i���V��bw���Lr�s-e�b�gN..jɊ�oa�����XL���OB䇋u��9�3Wm��T�/jX�#"⇶"����S��T��S_����_�-I�6�h	�A���Y�E�3��tj�
��{I�f/��[�9�!b`��52S�(.�x��E�]������+��c�mǦ �	�.�4=� �Ȗ��wC�Z�8��p����u`���$x�()*<֬��E������e�gխ� �Q�U ��E��ho�r	���$���f<��G�w�s��Hs		)�C|x�{�B=)x�djm� �UdO�;�RVV�(((`	QFQ���kğw�/v�)1�<<�***l���,ku��с�}U�����d����m~KK�M��Jvt�6��Q�&G"P��AeE%Y�����L�F#,zs�4i���d"?��DPt�	�i������ᶵ�p�w�W{�H���6�T,��U�^	�F����8M4��RVv����$�"�>�A�fbꮉ;5&��2�%�ɟh�/�Qt������B��J,pJ�����Vh*kAY���;w�4�W�z̸�11��:wu=�P����م��kޙ�.T��(i�`�ee�mnZh*Sh�˗/��070�'5-�$̼ ���r�W��L�O�hw������Խo7ww��z�T����V��F\Bc�"l6�D㓋��3sT�k}"����,��=Y��N��'�J�!w���������E���ݧ����Ѭ�"���.LE7l�<?T���k9}�8�>����{��L�;KB����,s�#��:��b�3%z6 ��̒�ig{������9�!�S�q����8$k1� F��=�������,�����v��]�����лM�.����f?���܌�*��`�$�!J��^�/3F�++��^�q�;���?^l���G���NY��xHHH�xj��VT��R� �8<,�~�EM$��f;�fh�������#��H�h��|���V*�(��E����ݳ�r!WhN�A�m�X:���j,'f��H��͇z��U/{TQ��bR���z��?y��seK�P��ʱ�W���W����zor�~�̔�ؕ[]N��������\O>����}��Ԥ}����ɩrAV]ϣp\�	��۫��o� b��=:��(:�+8�n�j��A��o(�*���%�Н��t����4�M7q ���)e�(��_~S�w��,�c�q���0�]O
�.�Mp>K~ܟf��$:���A���tX�,�:�|E�QRo��
ť��^�n�&d�� �D�k�=��Q��q�}&�&�XUL7-��J�x{��e�����(d�����6�E��|�2M1�����{���e��P@gW���C ��j�
/Y&�
8-�(h���ir��Azhn�:𲎛v�X�FI�'$�B4Π��%���a)�	<�rv���9��@eCl��ť�]�KM!�u�b2��/�G�Ƿ�����.�CYA�؅����9 07H3F�ҥ�?�E��LdP���Z��M�V�7kc��XX(�q�v�e�Y������ W`��&�	���^����.�\aEw. �	zh�K"�;K)�dј���f;�6�s��jrC�U�$����i��aS;,%������n�b-�=܍��6�E����O�KE��b���c�]���TP�p�qЫ�ws7+�_Ї�_Q�LQh���e *5��y�9��g)cx�`�.��N}�������G�/1�"�)
�,	� LK�<<d5`'���3�V�^�H*|���d�jyyy��~/ ݢR���z�C)lD���d�t��TCU�{����I�w�"���#)"�K˦��j����M��*��=4�K8������ґ���w%��]�X	Z1F<�fs-���*�F8?7�v?�:��(��b����|�I��׻mFWH��$~RiF<��Q�ׄ�l��]5��r�k��@ρ��| �����c\ˡ� '�ޒW����q��p�&�,o����J?����ʟ��Q`OG��y��O֤����L��Ӟf��n�l�F�u��5tӭ���<Tؖ��Ӥw�E|@�f�=��:[魤.,Yp[n�Q��/�f+v�lR�}~ LW���d��nYr s����4��붭�2�|W5'xR�����nh,$U~mn�]4�9�� �Y��+���?S���-��9p�O��Xvr�#����d StG��*4�P��bcck���~|l�����6���L�A��L��^%��}���I�w��ˀ��s��@��8���)r���>1��\��뮾+л�����>��kXN��\�)s��������< w�vE�I�O�O�aR�$�����A��c/Ċ'?|/��e�	~��L�=,����[\��;�G���;p�-N�e����V��(:���g7T:����w����0���h�C�������������W�"|��y���6]�@/�7�n�����Ծo�iəB��'�P���0(Vu�X[3"d6�}��D>򗧅&P���'��QІM���]u����}�S�K���z;�PPW�Y��}u�Ϝ4)UU<���uɘri�0"�{�{ڱ  ���
 ��fL�!�;C�k���{�K�>�&x6�5�rƿ3�ï��c�S3�DLﳖ}��ED�z4"*t���(ۯ��Fq-��n`�u�{�umE �JZ�En�L�6���D��{��'zM�����ZX2��A��v�P'�'<�,�Ѧx7;Y�����f��y�i�	�����u��8$5/��͕�+����N<ijokk�����5.4�N�9�)ݶ8��ٗz�8>[��=KK�-{j�א�F��Vנ�+	�_O����*���$a�.�~�W��=A>�gM�}(2��"g���q�i��(��i�������^\�wxw>I"i׌�]Ɯկ���C��D�+�5�v�:6��"��4�~3��fH�~_���D�YS���~c�����n��.�y������I!gU�Ivy��=���1����hCu9�Cn�6��� �Y����I�^��]�������j̊5-������?��븎QVc�=�z�x�<�h��(�AȢ��B	뷤�O�qcnGQ#/��gQ�gҨCM%-0M�z�!IsҼ&�ײ
	;�2 �N}`eg�2��BF@���Y��o��P����+�s
�$���d{Xr�rv�
�d�1Nt �F@�f��m���'�=
�S�<�?��F	�"1�n�����1&�Ox�)��.,t*t-?Ͼӟ�x����#��VV�I��u]�v��R�jK�8�K�N*JB�W��?�D^b�s�nrI'�����ᝃ��~�O�a�������-̋!�UЯҕ�,��U��v����mu�]�����8Si���2�"���K��U���ZV��%�	.� N��OMM��&��/�n� 99���9l��Bw)a__��z��ι4qګp s��,�ĄÝ��Bυ�s�yt"ܚ�J�乨$����A��͢n�w�����乁ŕ,�B,���Q� �E�H�����x��-�@��5YW�9�)w��ᦻ��
C׈��[����Uפȷ�q�ç�C4٩F�zxR
ʊ�ޕ@�:�<ʦ�2t��W�lO�_��x=lo�p���{e�[���0�p�ɾ!�s�5�&JeC�AE&-�z%� F��Ù8z�W��;J-��KK��3�G��J
�`�̱��A�*<?��t!����Z>�{}\2f7F��7(���	Q�e�u��Vsfu c̞�n1g��*	���O��^��bjL�cvN���n�-�80��B����_0YQ���ﭪ������߸����[�g��9~�k>9�u�r�y$bJp=���%��~Y$r{�7���y�W �Q�ZOU#AӢ���2>�B��Q��j�4$��e�w7)W�,ߒ2W͊��,DWf�W�Q���N)z� >�����
��.��n(w 1�c��y�.��\��eOE�]"�f"�Zv�����w��FDAÍnU_�������v9g ���w�����aNu�K�̥����"���K�K�~5R�#'m�Ū_����ب`����	r3�Ö6RZ[�\�Դ�K4^F��`��?M�4S�E��������-{n��#�݃�����8�P;G����g��
K�� ��P�/54b��S�~�YN�S�jj�Hq���|��yDE�$`t�� m;jJZ)dÿ���X!	,�9w���CA������r�|�a��.��qR9C\5t�>���v$�a���3����@˒9�(/���h��l$o���Ő��/e��Ly��5x�߀��c��������D��(^OW ���Ki:
�'��+܅�����pO�47���O+Y%��Fw�+
�3LQ��wS�i%Gʨ��4{���ЄoN��>�f;���Q��B��[k?���Qz��x���,����7�ïDP��]���M$��co�Bu�m�&`c��`�5����Á7H赮�M�=i�Ρ�y�x�%����A��Oo�0���v�Y�B����j�i�/��^jv�՗���̚�14>%��v�s��`�}b��Zk��*j��Kyp��~$@,��x����v�;��"�	�t��h|���T@cE�%�
U�e�f�*dύb�;^TTL�Nh�y�@/swjı�$�ߥ[5nv/��r������G<ﯝCNG�d���6»��]��Y�p����V�r���o��$=�|�6��W��t"O��~vV�^$g?��P�\l����xpEt�[�_���:�,��xc�,g�y�<�R�o�R���^��Q�oEFpc�3�b����_��� ~A�#̩3����ʑZ{|(Լ��}����
��$��>��G��c!�#VR��K��V������7N>u�%S�~:�����{!�Zo&p; (�gv�
.U��%����Ֆ�����`���w���y|�������������}����z,'��ɼJ#%;�7�W���k����]������eO+M��sjeP�GP�w�������7S�CPNUA��J;�
�E݋�b��|Ѯ
�ޅ�9���r�b͛V���)5�����r�SAXծ4K!�,��;��'�ʪ�H͘�=��a`
��خ�;J�[�U�($`�[�e��84Z��_�}p� �kw����oy?~��~9d|��b|��-:�x�|���/Fy��Y6{�|'"���c��eL� �<d�}����Z��M��o�e87^0?/.C-]X����\v�`��W����t�As��'϶`�����?���M��id����Dm��Jc���9���y=v�n��S��?��@
jc>%'C�����'��ScG�=rTc��-h�9��$X$���&��-V�����n��C�Τ��V�ڲ��R��ĎZ���E���z>��뼼��7o� O21��ӻ������~h���� �
�n���{�Bvt�T,�ی��b�h+R�T���4�]��aו.�������B�e3���T��ї�3hyI�{`���~u&܆X���u]U��7�#�K��)m��K=��	���~L� 7"���`䓭���C���i=��{}�_o�@핕����pA��l���[V��u_��'ȱ|Vi�L�A��[ O$O��*ѱda-'�w�n/��@�����f�ʵ�c������C���]�%k���I�f7�?�?�j�E}��O��H�3�\�>����|�Q��.1��@���8Ѭ��,8T�J����e �+8��a�(�K��jdÒ�������ñ��,�<.�$��r"E��}:a�}�-ޠw �0y~��\�{<)Z������I��s�{͸&��b�4+�uX�!S� $�8��IU��'w�0����zq���T�U�,\D��
}R����#��-��ˉ��Ȓ6m��S�$R����(�E'��n�f�tdQ��ݔ�5��>(����C1a�We��9;!���|"���o�֤��f��&�+��?_�@��)a��.Q�N�M���79�ol9��o��HD�&����2�Jq}u�N��B5Ԉ��Osh�j�%�r��1���J��|H���:�L�����g+[i��Df����c�*����ioll�x6�X!̷�ߏ$a�` 4Xj3\P�jZT&�C��jݿ}�JY2A�4�7���H��+����_�E}����<Z����o���]���E$�׸��us&y��&%��j�� �1�IJċE'���֞�����>̣�TK+i�� ���E5T�
P ����)������I
�U{1��s�;^�ԧr[�,@ls�����uELN�`�5�}��٧��B'f)��><A+��1C�?��tw�L�U��!d�]j3�t~
2��n��Ӱ0 ���`:Ō?����(<k%*�#4%^�2�l��2RM�i�G0����������'��?�"��(b�"��;�o����.��Ci�c%���8��<�m:�&�[����Җѯ�y"zzz�.¯)q�6� ���5J�G��똠��Z�י�d�t�����oE ���+�0������6\�|���i4S��d�чBa����q6BD��knSZ�����%�/F��h�.�^ǳ�z�cx��!��O�S��|b�B`���������it�"��[x�G�b�Fc��yu�Є$��^S*bHg^K$�%������%^��o�svP�<k��h �?p)���%���U�3~�s�2�K�C��y�28	�,{�N�kD<kG3�P��{kANчU�"�Cg�O@7l+�Y�>�xJ���\՞sM
�b���3��獭���薋��׫�4�#z���'�dq~�*e�2%%��jл�}A�� ��c�
���q��p-�ACC+}����T�_����R[(Q�e'�G� �u(d���n�����p6��-'�PO�Ȩ�0
QS��2!�'�B�S���~�kG���=�ʭ�#��OxƓ���W�]�_�W�:e�>t���amXA�˾/4�J{'���,|N�d�|�˹���K˕����&QC��%;O��^JU�?ST�$���ٶ<���Ͽ�']z��� jɗ�Y��&�TE;����_I}�ZR����,((QS���A�Pd�K@����W��wX����C��Kԅ��3�+*b쩰3e*�� ˩cf�z�=.��f��l��0�s�y���'��Xf��ot���М�>�p��h�`t�Z�W	��(SR&s����c�7��Ic�;�G`�uv\K�#mp�0Mp&�;J�c�C�]���V���@�W���\��x~�5Ѱve��&�5c�j�C϶5:�7�����T���ۚ;�r������Γ��k�R�U���E�����]�SԹ~�Em���y:c��"�m�U�EX����d��J���K�j���W܁P�g��g}0�AI���m>Nd	|�6��� ����B �2f�r����a���v��
�R`1�ʤU�O��K���߄�!���	Ʈ���D*�⪪�!�G;��*2�[
:)a�AKG \�g��$��U�~�M���|���c�~������"-$F����v��]��؂�uφs�|�㙹�Q��R�"�Z���A�SC�������yp"�"�1R�)PDS� �%��֎��FUړ{���C���ʞ[����D=@q	�d�s�J�A̅G�R��]�*{FHò��}wMb,��������g�s�����^��0�6�}�ΊG�M�NK ���YU��L-�r=�j���#��ss��>��u��}��!ѿ0.��]S��@ �mǈ��%���_���n��6�Ņ<�?�WL���o�s����a�хk��g�@�L���͌*����lj2d��Yޏ�8HCB9�@ՍՌ%�;�*����]$r2s�ֺ���o|`A'gJ�S�׾"�g^���&���{nz��[����]!Q��2�ԡ0�1�w��}K]��  ��������=��g�����.�;А"h�1v���yu�/J���ss�wփϧ���͍����?�����I�Ѡ2x��W
;??��a�9�_KNDs3��BQBv��N�!&!@6:2|b�"�*������e��3�d�+U�Tu:6��8��Г�������*��/@��F
J
�.����d�^x�Y��t<}����Y{�� ��Vƒ&W�mUӸ=C�	�5]a _�!���n�-��+I
�n����/���S�DCz^=1LVu�w=�O!M��u�]�k�U��EgT%Ɗ�$(?����&�	z���у��􌼝#����'�����n�bl���E�}�-�+B�p ��	B�E��KI=�&Lss��}��pV@ �ïu���l���t>���������
��^�������{*�r�aEE�xLsC�����,�+"L����s����:����B��)˰���	Z2����P�/nD�S{��ӈk��6��������Ձ�(s�%/�����R���#���:���Բ���\�ڊ^5��!���K���j?Q���9B��qؽ��s���ZO��t+������}��<�n^��䀛%j�2,�mXk��0�^�ᑐ��_="��������?���!s,|���Lp�0i
oI&�r��t���5�ѬG�o�~�|�G�qM���T�����3����U �\�]�V��=����QǣJ�O^�Ъ�B�4a,���7�P_�Y\\���c��<OI�bY�J��d��u��5:��Z;���a�L̓�������I{s�w��8P:o���X�(]��@��y,(�7 �u(
�^��o���'� �
�4���t����ht"�T�N.�N�>�Xd���������6~���{�@�&j���yz�CU�/�ޗԗm'TB��U8��#�V��j�E��[�AO�ۥ��ZF�Y���)5�� ��ȱ�p+��uAS/���o�c}��&)�����Z�D�� �t���64h��B� >>��矵��~�b��073��q��G��6��4y������R��Xl�ps3���Ⱥ��L��-R1��H���H��������ё�%�}�'7�8�9	d��E���^3��'"y�TTTNR�p�y#q.G��O!��tS�7���5JN����O!��zNlywN�:V3j� ��R�,7B�C�{l�!���S�g>����4$�:�%*��FZ|똪�WˉQJ���$c!*r�Ӓ z�pۓZu�ǳ�D̐<ƨ���C���l~$��(s����Z@�o����6�|�)�WR����"�I2�_��:޻_h����Ӥ��,�˞/���X�����5Rq�uww��>^�~���(���$�Hyzzj�PA���H��j�Qt�X���||E͸X������]3�!7����
R�"7/oXIII�S�K)2
��B����h�ǖ)�ᎫU���=��\�3/II���H k ��-礬��H���@�n�T&�aV�E�s�p<���3eR���{gNX$��.��|775���Hc�m��2%�tCp�˼�]�{����:8��KY\��xCLR�+������|w"�}��j�-�M�^���E�� Hrz�*���/o��ʴ�E��LML@�շ|A����c�	����/䍶������L/f7,ifu�;_�@ߋ�f��J�Q����֧K�utuK}��6���|KK�o���p�Fr��Y��nncSl������!&�i���eUU�&�(��#p^�5� #�h!�W�h/G�nx�Q���^A���#b�y�o޾����3|�ƚ�YF�p��v]:���F�ɶEo��C�gF�#�&/����8و\��X ��F�GT�ʫ� �w7���ѓowP�U������+���1=7���.�E������1��������D ��-���leCC�ť��}�Y&����<���Ԙ�11�\\��S�f2�
DX���c�J��FτF����㱥pK�?�����r}�
7�����#JѲ{��P�F�NGu���ޝ0|����R[�R�c;��+W9���'r+s�=����_l��ϟBM�]�������(�J��PYA"����*>q�k%�Ĕ��`�E�E���RO�>:��1�X�4��O*�D��� ^v�*v�0dx�A}�]Eu�Ǻ�e���o�z0�i����W�6�@]v�v�y���G+GFU��o�̹��J���mHO�TG���6��ϷL�������@ѱ��d#��F�51q��&�̓��`w�d^@�	��6��c����v?����r�k++f�%a���J'��=���[.��4 �'�� 1�sPгP�ܨ��C���]>E�e��Hx�ϔ��Ņ�gu���f�=�v!����~��v�6��K4z�w�t�Q�&
V�o�7qr���y�㲑����U �S�s���5�A������֕f�=J�yF�f���QV� ���p�/a����v�j��oٞ�M�r�R؏۩�^tR�j�2����:�����z4��j�������L3�Lp& Et����9���8h|+�=������p����᮸�54t��% �h�/$$d�����+�`����H��wh��5�^�l/�L8Mf+�����҈�/×�{/t{{�)$T���ڤ�:b�x���̓/��`�=��_\ �L�9�>���������yxx���t&�b�Yb"�*^�	; ���e}*��S�6���A��gi��,�����*��^ F��9��	�d7���������ep��`b���jlg�#�c>�c	7a �l�8C�VՑ��~��#D�+���T��-~F����϶{��UB(�s]�?��3�y��%7�P(��*z����������1Q��K4�mu	�]غ["σ@E�Ԋr+���K��jGGiF�Ro�;�Z]��Q�4�Ҽ=�+����"� ����MZ��^��C����1g9Y y��# z+�`b�_�up k � �,V�����8���~4T�J4 C����mw�o�a�o���ohk�8��D(b&���J���?��,���"��D���	L �Bu��٥ S%�A��@6��H)�h�3���ѭ��L�2�V�G�&��~���z4?�}l��s#0H:��or7`�w�u�z����M��)*��)��p��������gC�����7c�'Q��4l)g��ns������ +��~���}ÇI�B�����?gR����V�a�t,��E��S
P��~i�����6�p2A����]�G��4�I��W��7�ij�W�^�)eP!��kY�������������1n�;��o���� ̃�z��$ �`^������	ۅ	3B�b`�̙��i#�Jm;�f(��Oҵ�qF	s��L�k��9�~hfy�<�F�>g�ֶk:��Ͽp���L��<a�Y����{ ����;F2^�pPDʲv��G~����(�eQ�H�o�Ao���BWy�� ���h�q�Gc���##����؋�L��c��*��ĹJH�������/��r|Ts����.����ވ4fQ���G.�v��t�0�g���3�#���y�kuC�
���z͈������Z!4Y3M�2��_�_qd㤸2i���^�xP���Ǆ��4��*/,;h�X�(�������ZBK{{�.���&]kaʫ򫙐�����_jd��&#5?(a�zj�U?l�V��S�3W�B�ӼH?�c|
��rH����`�m�w�agp�[@��uJ���û��4�]�'�P���G9���'�{�v	0���lh��s��O�#x!�g��տ��`\�7��
o*d�ʪZ��KO'�L	h����EbhnN��Pҿ�C��ʚ��Z��111��<<<ŏ�o����3�J�� �.��?�4��2��,�v6�|�����W;]�ѿj7��6>'��(7��)1I�}����1!�'OR��k������g<�������Sg ��G��-H_<�P��u��*�W��s���.;;��>ŕ������I��X�|l;N��p?����f�.ƃ�3q#�[�:��٣�		��F΄D��vǕX�m�����O�M�t�������l�jBs3x��^ޕ�&�&�f�*�_0�ϦD#�Q^mF��Yo��0�{�N7�����{�o�5eD��]��],����V�z*� ���ߨS�d�	�O���M藭��w�~�b���2�3�ېΉ������4W�^m�����i��֘��e�9�8�b��y �h���j^}���W�cN�nO��ud��Y���1��[ck���'s�:C�~�c�aNcn2wڗ�&�L�f��RJTͲ�����,?�l~$�x�3�!R��>L���|ښ>�t�.ѓ�i����n�8zNd�}G�<�bꯤ�F�=�B�\�8�ZŔ^�C�S����T9�
@~��3�!�̩n�5���Κ���3"Tc�ģ���:0�Fj�Tڨ�F����T�c�dk��(�C�F��x�*�߱-�	郞^#�<(�D�1�@�˅N^K�?�Ee}ˁ{��%Iz��^��q��}҇:�9Ra��� jL�[���.M<u!q����'M�M5V@��k�m
]�͘6�#	����t��N�'��X���i�)y�2+���#q tW�v��� }CZ��6��9���ۆ8{�\Q��3�����3���ֵ��)a�,�˛Q�^����������zg�g/r�C��ڡ>�:��5d[>S6�q��|�-ƛ��Cs��&��-L�r���;~=/m^e��M�>Q��4^�
�4�h"Ez-KA�Uf�$�-$��\D�dG�t|�+]S,�U�Y�?��d�	��T�U�\X�V��,P����l:���qZ*M�V�&4�;��tpH/��Hߊ�a�Il�ܜFڥ�e�T��5���Ʃv6��� �\J�M�M������G��^vUf�����lfokN���d�ES}z���ߜ�@B�s0U���GP�Qn7�{'�늳��	1��J��x0��>�;����)S[m�����,��q��5k�<��ZM�J9�ޖ�i�`~�\$��,���՛��=ܔ��5TGc�{~�7�������S��{�C�`y1�u��H�`����d�0Ҭc��V7w���o{��E_y�P�}5�?}��w��GV�s�R��\b`���W2R����F�n��b������M���J�l�(o� �w�t��%>锕�p �7��e�h G��_�p�[�;X��/����?�׿�������H��IӬ�_�[^�(]]\��*0k��ءw�Լ(�7H��薘JޗV���&c$�uCa�Κ�����w�*�%��ȖjD���=_���o]�r`��C݊��8��1��&����:�Xz;S�u-ΰ�J�������������h� ��}��q+�W����v[�%���X�.��P��8k���֟��_�W�
s+��(R�OX��
��'WO�φ�^U\�l<����ox����B�$B���c!��$7y\ �T�ͯ�ͱ�f	�݀��ñ��v�u��'�dM�@d S��cg5�Д!N����}I'D�Vxyц����f,�1|_��m���+I<.��).���q"]��%� ��1�� ��RiӶ�Sf�����H�
Hr�}��̫svt�6�SC��f'�mG���Q��)9CP�K8��9�A=~��2Z���}	�k���M�_����m�^`m��F��O4�BOte�����TY|�_!���k��?J�z�`��y�7�;ئ��V	$ .k,3U���b��T�Z?�F(E�"h��
��)Y�3���Bt�-Xv�X� ��#=����=�ۿ64��g�f��*����*�S�`mKG48���V��
�%�6�+9bQҗ4#)m��+�����?�ݭ\�4�u�՟􋱣{>'��үd-|V��^���I嘣N8���4iz��i4�L��
o��+���s���<���͈_YI���ཱྀ�DsֹT�s?��&����A.������C��?���
)]d#?�J>7c���?ݰ��D��{��>n�q�pW��B/�$���p�+�we�x���V�!>����ꕓ>��,]�P.��](����4�f0@N.+�o���^ƺ�s��TŃ�h�Nٮɂ����Pz���(7"d����r�r��$����¶�9����uXn����ļ�T�v���X;��?G�2,1%�~��8�[�5?)2����y�^�i�h�<�T��;�x�������!�:�r�L[h��.S��Akc�Y�7�[���g���q�/MيD�A+�:yN����*����	�_>���z��ǟ�����yf�4�:,{���1k�`���R�����=������Q��֒�)�(���|x�i3���Y���حj0�,(���y��܃��*O�L �Wjo�����4���iZGa�&��y� �i�,}�K	���	o���|pt����[�(@����xٻ쇯)s�8u| ��/�:��=7�åWS��)�NR�?y���Rg�{>v���@z�x!�Ђ��̫�ܫ�+��+��F�!�/1��;��3�c�k�$��$�x�]��M��ׁ�7J�䃑3׭��v״`O �Q8]�.�P�_!�&s�ԩ�J�E����� �n���2be�I$�JpK\�^a�oVr�*�!�Cr;ޘ�Ǯ��;�߿fl�c\�a����Z�d�5�~���6���`���y��5�N���M��ǿ�a�7��w���b6�s��;��|���f
,����;4f*�; 7I�Ė8`So������iRت|�|�λg;��ʆ�#iF<����1�\||�K��Ģ�x�>�}^�6��,�����^w�b�u^]����&�k.V����br���S���h�T���ea��W��c���~�6���K��6bI��?�*��C}�m�F��@�1��xI��u;a.MA�ֲ�G�ZG*fD��X�|x�xA����2'z�QS��V��b�z�����i�k�/fSb7���������o��'n�����hԘ��k��ʚhuy��Ⱥ���|>3F�Ў�+m��۰{6N��﬉�vK2:;�t�����-E�]���l���^9�rȑ�,���3�8���Rp���р ��(����'�oö#n7'���+��l�گ- ��
�CF8_�\���ԏ��|zI��Dz{wG�Q�J�������i�݊�����b"l�p�B�R���j]�|�r���)��ӗ|ъ{�e��S��վ�����I�ܳm(�N�ү�e-��O�y���=%BO ��`�ç@�`zO���,F����J�O�����=��?���R_�_�#{o᪙��;
�C�����ڎ���[y$d�eee�x������}#��9ͭ4��UMo��#��q�s������D�9+np��('�V�ԡ=�/�t�pZVV�O�O������BdKȞ�%3�\{d˸�^!;���̸v\���������ǵ����������%�s>�y���~���A���Fi�Q�6\�[7����q�5WT��̒h-kd)�K^]H���;+�%�p�uk�'���u�;-=cŰ���z��JCע����*�:�E+8���M�R{m�h��ps�S5E�AcH�ᩘ6��L������9��u��Z�{ē��:�Nܸ�<Ct���Mm
�걓�)U��\��^Q�"�k6�)��*~�y%>R�h2bo��3�U%�9Kx�~��G�"y``l��vrof\5[\�)�����]?$��VL�ϛe֌N��,�,��soJ_����~�=�����tq,bZqNv�ܔ�����mQ1R�o4đANi8^Q��Y�36�#�_]__W�b�`���̖��N���׊��H�J�2k��ž=�u/T6������H�7�6��{ec7~Jo��D��Eӄh���o�Q�U{r�X��g���j�g���:xp9���!���*�1�ej #��,�r�L��rI1�~�`�z��OV䘣b�ph.��C�����i:Ў�9f���C�q7�3�}���E��L�<�I�W��j[�4~��/���)7�6o�@�g���kHq�Lǃ����������e���	[���V���Ѯ�.��\�͙��३��1{�'�d#c��{ag,k��D��a�t�N��j���-x7����F���7����s�w���3$|Z`��)�B{�g-��j�l�⶜ud�:�H��:��o��M@�6�BLl߬ꖄG�2z����\7_�j�n��C`�Vn/����Dx�͹���ī�w���\ z����1:��jl�G�o:���DU���{4��`�&G�%�sl��_�B)�IV<�6ǯ����+�����0�2��A2@M/wϬ�o�~�=�rDb�s*x���ks���]����?G������V(�q�_��� R_�bx�j��A�P��J�.��	�&��'xZ���un���ٹ�d`	I�����6��0�S!�z�W���%�L��ɚ��$>��9��E�����g7�s�N��_
�?��40�Kp���eXNe��|��}ם�K��1�欖��ˁ����ee<��7���tX����ҁ��/�D8�655�D�����gc(2���`��6{D�i�m�=ߣ�¯C�ɷ���;{�ИRƀ�Ƨ�--��Ҙ;��B䰞={��CK����C~j+l W���c��/��t�zzs{���"��K� bԮ�em�.2,�
����OW��:CF���4]Pp����!EG�m�91����H�\�ْoۧ�Q
�?����<蹧r����8���"��y_眄��F��[�|��$#�n�8�B��9����5խ�k�<|��C�"�Z�.V�Zǫ
y/s9�`�z�)�nȽ�e��]�g��Z"�S�jl$L���J\�7�}�n�-����3i�sP�����3�c^  Ռ����YzzR�鸿��O�ĭ�}����8n'�Խ��K|?�yxx�śP�]sp��ɉ�cm�U��^y~�W݋��mv��/�qr����_�$C@V6A�2�o����2���;Ϙ�T*�V0|���b�n;�5�Aw�O�ej9Zr�L-��rي'�\$S���~u7�yW뾼V�H�Z+�v^*�Q��_k��s�^D p@C0�܂��h
�y?5P�W���8�_�)���� ��	pu�ݮt��_�l)U�[�r8T���ڠ����Y�ni������'��Y��������c)����x�{8uaԯ��љ%Hư�h�>������?)S0��0�{��X�Y��4����a��~�!��j���0/����ׯ�)������9<��ӿ$y�2�24��h��I�v�?�L�����|m��u��x\�9<��)jo_�	��J�{1���/K�6��`�d�ߜilj�u>���v���?��E����[����(�p�d`�K��R��e\\\�Ґ�
DD�a��^��-0���VޔM@����{�{�P&PD��`.�]�7Ͳ��q��O@��p��e�� 6��H�Zn���q F/E�:G�s?�]���OT����J��������l��g��E���{��.|xU.�?o`Y��)g�p]�6�u�|��V����}��M[��g���\���A�sw�������f������{�n��"��wYY-'��:Z�ȰNu2����&6�\�yӪ��^+k1:En*Z��W��/Lw��ܹXXU񦅡h<W������2TiEE��^�9f�v�_��Oo ��Vx;��RI�����M]Z�䈩w_�}4��`�K�ҘW�pi3��1�?W4����6�M��9����K���n�! �2�~vS�2ޢ��b�fr��Y@��>�� ��ӵ}>%�1�F�-�?�((���e&̬|q���
�T����Z�3���=i�V7��m�e|�J�iP�{�S��×Lj�R B8Һ�}���`��AA�J	4�7q���tl�� P�i�3�R�]�M�qy�L����D{GG�r��������B�~��1" 7��n�'Q �:Bn�ڥd611�SFx�g��W�-�Z��ơ �}���"I�4(J$?�<	ֿ�y<���2!���J/�Hc�Q�C�Մ�J5A֤�6M����3c	��V�_6�y�Q��1;�BߧĆP�;/��F�r�.K2bA4�R�5#-.�Yȓ?63�m=�etF0�P��JP�n������C�$SM�>7����_��
<"!����B@�	g��\�Ѷ�A"��RF?��V��rq����(�M5M.K����Zv[�$Ƽ#?�wV$�hW/�������N��-�M��w����L�T�
���LDB��W������ZxDEE�π<@$��Ҍd�}Zܶ�vp���Z�0�dx��j6Xoe��D�|*�fɗUЀ��Լs��$*����d�7`�ڎ��#�U�eғؗ�����K��'�����O�h���1c�����	Θ�sd`/��Hˡȇ�̩�����E�����x��1 U���,�F�h䀄EA(&&ֶ�� ��#z��� !�������zht̂�����J��5�vnoHy���x��ay�`��]_/�n��@�C2�?a��;�n���j
��j4�]8:�VRR����Bypp�˝�Ӧ�.�yg|��[��7h ׽N��cr�25,��;��(��H"q��n���[�ӹ�4UL�4��Y{�0��-*cʛ���&��˲n���[Kʦ��5K��k���8Y��,I��G�We������/�)sѢ�{�@[1T�ϧ�9��P}�yi؊h0���q��4�Ud�?;���;��75ٔ��i�������+�}�;�!��H���0�����<*x�w�
w7��2[����c�t�r���߿�x$�JX���Q �C"�Б��&s�
�v1I��/_����4603�ecrpo0� ��o�`�ȒX"�׷���c(���}`C:�!ښ�޾>
B�W�|�lط_v���F>f	1,ÃB�����:A2����E��Ӊ����g� 0�,nB��It�p��xJxyy%O%��3m
!9�C�ףS��J�J��1���-�>;0�<r?��k��uoOH6���V��I�+�,zF����a���>�Y�f�gGcy�c'&�khf��q���D����׉
��|GYl����]G����gd�.�ǭ�����UO�t5��(��ObZ��K���v� �c5=�9�f]�P8 C�=���1�P��)��7�<B �Abzm0d��9��:��,:x���Z�E�|�t�Py���@��ǀ7����kic��en�mQuu�h�c�L���(��L������p�ͽ��1=+�a-��<J1\����)H���kƺKu���#���Gh�吱���2���)�v��@g�ͽ�7�=���Z/N9�C$�sҿ\��G�`+;��V��=i%�wI����dt�n:��7�*X*����_��7[gH�&��l�K�i8��)=#cП�������^V
�)����u �a�%�1.b�1�Z~l݂�)��)1��4��mح_v�*/--��G�ǳ�D����m�%�ǂ�y�,�:�A���Ւ���!�� #c�a��{,m(�1CN�n�O������%h��ҟ��L���X���N'��>����mҋ����o&>��+<ٷ'l�Zܕ�P��������X�W:����_��rG�6n�'�m+���2�YY6��>�nt�Q�I
,�6����K���u7R���V9�����F��^�鹉�+��L����3���2)Ɇ~]�ƹ,V��e�L�1�����̤?~av��y�ix������Q�
!�u!��M�^;�E?�gx��Z�O友�I����*&20_F\t$B#3�_�WnQQ[�5!6i����\�ݒ�K������T!eJjO��-�����bb_�q��@Z�+����8\[�4$�~����=yI�+��?�Ɯ�Uu|���Ȉ޹�}oa�s^j"{��d��&.��)�O)�|�y��Ƶ�o�+���k�޼&gňû�x9&~.��2�ɱ���K�����\F �xҢ���ND�..>�;��8v!�^���n�{����5��qk��������Tވ���34��l$I��n�k�W�@��L��G�B�|罚* ����䚇��/�
������r�OkX���4�����~~�ͧ���Փ'k���MA�wfϢ�i�����
�ؔ����I��xE��U6��^�M�꯻%���A��9brW|�|Ŭfe����f�n���Hf���dؾ͆r���`���Ms����}�[�d5y�W�6��ݥ�A�"���(.�.�Ə��?���]�ڡ�x��p������N/��5�/����)�&�{I?�}Kst��}�p�{�����
s�6��Ԝo�����r�<��sE��;7�y^4���Y.)U��qa�%1>$a�h 2De���<����<3�~e��`?�k=�<��� !��JW�[�w���LD"�UB��1ǢZ��(ڻ7C?��`��Z�*�U'��Z�KO)'��fY	F?���2
���s���*��G����(l�|��6}��
p/B5;���i^#�<�~���_��#Ƶ��BG&�%iT���tEd��Ӧ(>2b��1@#���c�k�,j�E���������:���yy�*s���	��☂��d)y�.4��O*��r�Pʞ/�K�u��0��aH�� rZ����I��3�7"�����P��Yq�3UD�I���ל�	Цk�9�ӸE���;/�T"��3�yB��FM �/l n|�d/�C'A��N?���s&����n���i��K��KF|���U��e)��=��1}�ﮄ�+�"1PP�z5��ÿ�MRCN�4~����GF~��F9�( }�F��b�,����o��uU�i�3a���F�O�y�DԄw2��#U�W�0�����Bv��ˌ�g'�E�\Ti>,s0R��;M�|��.6�� �6���F���Yӵ��z�'�#�k�V�c�,V�/��~l<\"`���!��%*�
3�u��P86J����m9]F��������|�q�0��^ੈ�嘦\��`�����[ԋ���9��R��C�o�Bf�K&�y4�`m��(Z�pZG�|F)hS��~D-���$��"��ZT�8�a\w%>��7E������#�p�>�!�PR;�sHK�K��o��du�[�GW�|���z$���͙iƼuE�:m���W��IN����W���l:�eW���ֿd|�t�+������J9��b�6�zZ���*9M�'��iU/=�(�g��ɄV�颶�܋�ae�{���ك���^˴�t��
U}��vYVE:��٤�Nv�t6�,��p�	'���7�]O�|���$���ˉ7�L�g�<<�v\3z�G5�{�U���u��tc�i���-��|���C�s �����堗U(86��w!-F�"�9��x�I!W�R}�-��a���@��i!3Zom4Ib�m��緷+���%�(b�'��\�c�J��'��~yڳwp^u{8�֚&EUa�|�PY�M�@ߚ�g���!�"9@f�U�:��Nj�E3�ɱ�<�l�Ԇ{l��W����k�t�/L�!"�z_ݼ�ɸ#V���7���*ID��b8g&��!�g���	=�P�q��6�no ��i��7�87�nR�j�N]U]~$�ϔ��6�^n2�bR�7�Q��P�Mh[@���~c	ܾhG#�R�&���*�xC�Z���g2�x̨�7em ����hD�%$$��}(f��z���&8�J�_�Nq�֘]�e�[��MC�R��`#���+9t���L+h�^`#U�T ��_6�%�B��ƹb,�T�U������S;����U*(V���ڎ�
-K���Oя�鰾��?:�Z�"���>BZK���r9p��Q(��L!|U��ax�����bѼ��E�u� ��П���GAx��s�t��&� #&?f�A�)h[C@h�u,PM��R�v`�p�Ty~���ja��3]e���~i�ֽה%27}Y�wA�������5�6�=��r� n�Ht%%%�5�X؉.S�VIzgF����̝��/;��k��B��m�$b=o�C�\0]ˬy}A&8�ף�e?h��+{�p>J�3�hq#=��>A�F�����1��^�L��\@���M����`j���쌞n_�:�1����7��#�0_�u_���Eo� _H���	=?e�Z�sc�ai6��������������Z�pT��ҟ�����)�q7�M+���9 Ť����E�B)e�S.��@26V�^��΍o�#�]���tԭ�����ER�Emr�����Y+z*K1�>r3=�\������WYf� |��61�E����W���1aF���7�"`ֽ$�M���?�Y@�
C�*��9Zr2ٌʈN��K{�~H?�E��q�
�eM ��C�<ΎuK��^?-~e�keߵ�`	��U�����._6�������|����^�^
�����^*�$m�Xrss/K�]RN�z���b�6Eg�3F�t��1e�.$)���Ϻ�O�-����`*��E���L�h8�
GZ��H�Mu�n��:]� �t�z�}/�����Y��h�ĄF����d�Q��ʐ��̏��)x����r����+]�s������%:��}��+++%-�J�t7��.�Oՠj�I���_O�0�>c�ȡ����[��&NJ1@�ۜ>�KLGG�����#u���ȣ�d�½���ޞ�r=wvF��j���1Kb=!���:��m ��������96s[���K�Q.�!������p"@�//ڸ#��y�LI���>=���-�q��b�`��&v����e��C8�͉jeo4���!��K��:;���5�4���v�i�G.����������>�~t�ga��s݂��g��K2�MU�^-�s2/`U9�Mk��f����ꈕ`���ǫ��W�rB����n��aI$p��v-
&C�@F<-f�&�z�M$(��;�!ylGeMnZ�����pn�_D亂��2��a�J�2�1~_j�������k�kcc����X�}#�ݥ�d�<x�y����a2 �=���=����2<��5��;>d$�_�������]=��iП�U�D������b�ĺ�j��O1�a���צ�ji)_9�S&8����N*�u�g�q�Ɯ�)�.�hB{v!eO�:��\��W}K{8N�ETC�f������_�(�����_o�5�>������ ��/��_|stx��z�, <���ḏ�'O����af����eрoef�O����sS�����eJ�K� �g{��ߥ��wL���*�	K�[����?��-r�k�mlmO�oW3���~�0������[��Ѝ'6Q�%1www�y_~��7�c���6}�����`�Ϩ>RY�#2�c�GGޥ�u�4��:*���8Pgv/V65��x+�P΁x�&zT��]jK�@!���{��B;..dn�lV��A ���z�]o�M�֌�ݕ=��,���'e��[�a6���0�A]//�[���.����`f��M8@���o������������ˉ�/G�"(((�?oxe���k�����!��zC�0Ϣz��i�8o Q�T�.>>�`ii�}E�A�h���p?�zkǭLGH�!��Z��Z�&�SG�xRE��E�ו!\�uoRTߘێ!<���;��� �IѴ/yբ�̵���U�aC�˓�D�X�$�M�ffl̯-�i',�Jv��?����8���k��u�!�i�wiE4w��Ԕ���3>c^��[ �Oϯ*W���ӦE�5��'�� ���x�ڽZgr���-@$�c�쏒X�� ��Z�ڬ�L8�ݒr=%��1KbU�`�.� ���܉U�1,�r��Q�Um��>ז)�����r/�wZ�ΉYv=o�?��Q,x��j�z����VVsN|��{�~���Ӧ���дZby_h�id�~H�V��Yh�q8�:��&�fw������͹��_��E8�Gʾ"�i�R]�h����׹J�~��idl$)������C�" P��Q�*�����/xW�&6�ݗ�a�]�a� �)���7޺C�%�mgG�=�٥A��*v��|�#dD����s�������ܐ]x���;u�\���{R���bry����+�1���[*@��u������R�*�ol��.y5UUU	�:��%?����|n�^WJ��	���6l !��%$�=�c��a}�(��!<iO��'���)���� ��gY�f9h�_~�����n���$��d�Ǚtk��_J��-������<�k���4�*��6�s��|N7�җ��򽴨��ؑL�V�&K@a*9VQ�C0���i*��{�j�$'H` �\�+�*Y���*��ڻ�g��k0"�-�γy�O�H�F�>>8�Ą�D��_�~���\� \-�h����R7�@�8:;�Iį��n>�m��ݛ���.&))ϒ�|WH����"�l�ð�Ƒķ�^oZ�;Bt��zS�|[ȩ���CƧd��L��/�]���)�׃�E�ȉ�����;�'_Y���	N5�a�Pai�C�gMS��j�墡Oo���5k�)�0ݍ[�&�J�*))NaË��p�æ�����!�Gd
ژ2��T���e2HM��Nc�v�1�eeh��A;�J$��b�+a݄t�BVf&s�� z��6�5��~�8m���������w�4y��Xo}��[�>.�{��ϯk�q{2��9����nu�;TT.��NL)�����#k�=AdI�3sk�u�$ �L���t�vvb{�l)E�_�Z¿9��0j�M(���Y*!�6�|�
��$�0��9��/�R�o ���^X����z��������r��zJt+sF/x(z?�4�wU�j[�R@#<��Q�]�x!|�̷���_� �(t�6潗���_77�CjA�}�lF[X��*�dGv/>���ڒ�I��9`X�x��"9����T�O�a��pTW硵ʇM��E�b�E����@i��@*�l2j{sݴ⎐�P1 �⠊�iA�#�Լ?d����(祇D�#�{2�A?�	�ٳ��������ZfU�Ué��A�|���:Gg��>�aH���D����r_D��v�w2���#�щ���M�z?6]�E�`������'��������_Q|+�m���T�nA=}}����o���}���@���0`�>|�k6戇rNY�{��^�~�B�� {W<XnE/K�^���� &4�H�@� �1:��@ʿ���mO�'K�j^�nI��G�*���jY//������{�d�o:����(���aG�1�G�ْo��ʥZg������gfu�I���z�l̨sS��U��y��T�����>u��$��Mu#��"s9����n{��+�*A�fi�����}�3Ѧ`�u�����r��^,�Ҫn�?���妠������G%
�������f;�T������<K}�H��Q��豩.���+�=��,5������C34�Ή������˟C �Z�(�.� �B�1��ʰ=�0��Py-��>�
E��1;O`�=k5z"��+A��W��� O�Iw�q�/6�&2R�C��a���ʓG���޳���[mSsr3�'�����ہ����eK����j����b[��n#�n|�v��JMD�{# �|���S�����N�u�u����)��ć(��1��J�r���Đ9v#d���ދqI��f��� �=x��[E��8K�v|�����n>%޲�!�|8�����!q
0D~�t�q�&\��k=͠��!�Ƴ��Ȇ֌����ѝ�qR�'	3$x��"��&���yH�oQ6����eӘ	�|v�'4?��i*�9��������>��/<95�\���~����X�v���f���}�zM���φ�	k1Z���)@�!�N/w�dBc��N�_����{��uٟa����l�P16�H��^�C����<��q?��K���vߒ�իJ�����h�@:�wh;��h�L��.�����N�Q���:�L��i�$V�ij�hVf�\�o�\Jk�b�(��y���KӀ5�-�ނ�����"~�E�.�����s2��
����7��A�"#��0e��y��m֧�Ȱ�]�Kщ�%Tk��V#�Ahd���I"�,?N�#��h�0F��߭�tƊ>Zc<c2��Ed�^`�u��'&X�;<�$����6�M�}bw*��eHSjP�������OGI�����*WH�\)�V��p���v��:�R��2n�_秕n�[�u[���P�`�#z�?������Ե%R	e�3_���{�Fj����e���95�vb���r� ރ[�c��u�?!
^���OEex��P�Q��MS~�9|�i��ӭ��-��sQ��vaS;B�}{������Ro4g�j|�mSm�e����j�i+r����o��
�_�:G1�H�w�$���ݲ6�p��UW�٤{��v�h�*8��OW���\�Pe�F}ÊB�!�td�C�E���݆Fz~ӣ/�t4>M��C���8CV�hd�E��+לl���%y��K(5:}�#������҆_�N�s���F�1A��Xڛ�4DO(�Q��6g�}�K��g�WNO���~w�j:������d�P�;u��ϯ9�Ĝ�<�62�T�Hsp �op���d�����1��u��Vi"��s����ɖ��̀5Q2���/#AG퍵r��ɤw�m!�Yن�,`��$�<T��\��b*ϭ���B=�_'���#�w�'���4�JK������~�F����:>�A|uI��ܿ�ev���.V�����g�m'�0Kj�2Ù��ߎ���Jȋi-G/�MCH���.r�"�h�̖���lg�J�6s��Ú�����7���UY@A��@zLWS���B�e�m�|�u�WL��^3�^l�>�&��ё��+5}1�?�7B?�&����%^<���ڞD���mt+v�ԝ/���\"�����a��S�����4U���-'_����A8����hD�e���d_�>��kCH���FA���~���G�����B[�Å53��z8+�^�t7>�hM3��RT���}�✲y'��DT�θ3��rHK޻���w�����fÁ-g�7�~�n�\����`�ڃ�?�)��Lc�)�pl�Dv�8L�Fn$��rCjE�uf��B��/xF�
e�:��]�'�|�|�I
P��/=Q�4U'���C
}��Q7>{)�*Y�@�oe����\��O���G�g�4K>���A֒G��4r3g§�nL�K��U^�d��:��j�W�۾DU4Q���R��������=��%������Bh�H0EN�b������+A�K宨����i�wS��Fa���,ߊ���͎�7�{-|��,�]*��ԍ��J�Z�'v��o3��!����~�
Q���H�����`�ʄhR�-�����_:��X�*1�s~���yOt��:����#��(G����}�[Ђ�t�+4�D��������7Eկ׼�6���Q�.`�'he����V�yZκ���)���v&i��H��X�a�|�Tsi=c�A��8ɿ�L�UN��N�\@����������,�
FB1U�IN��7��;"�����R��~�����i�<l�s�gwyR����c��QDkv��}��(��G��〵��0��.�TV�v��0>�*s�` �KA6)��.i�Ņr�X���I��r�.B�
�����i��'Âm˞�qs�>[T�W�.x
�yRBQR��!����E�g\o��qfr֢�p���^<"CN��1!	ػ=��p��M��m�_��P�>\f����vO�y����|�U��5�ڏ�=?�9�ܽWϊu�<��-��^X����Ss��6�_���q#'�{�nf�qD�k������[�&˗�R4��\bͷ7�'r$�1�4#�X�1��]<,,���� -����܃l(T�1�0�E7���K'k��_�7�u[�C�h���ZK�%>���d��|{���_��b�\�F���*Ҕe���z4A����{���~�$흘E�rx7rA�H�T��*�֞<�
�J���\9"��U�>�.	�'ș�)�oο�?,�T�rz��{���xY�U֏ϥ�qi^�rD���TC@ԁxzƥ�4�X3_q����\k��2~�C������� �����SYW�]k�ß�˟�xY�;��������V���ޚ�Ǝ�10����yF/��M	�g��@����vr���+`��u��ʬ����t�jX<br9I����[Q&K`(�ק������7��\իb�b�
��p lh���E�"��y�n����i�����	��w�c�L�WkS��w{D���z�AO���=w�����	����{�}Y���+��M(���ѵM�CK�%h�����:f:{�)��n���Ԇ��D��H����E��<)btJ���~���J@����������F`�E���%�����J0�긒Aꀝ�Vňv��Q�W9(������I}+ǸİLJ>7�A��F���1f�6�?W�V��`v�p
ܖ�23s8H:���&�No��4�1�u/IG��0���aX4la�q���L����8\�4&w��7�)"����9�U!�#�Y�������a1@��*������"��{��I�h�ɢ����D�+"�V��Ѡ8�BM��H^�|-�r}�ģ¥n�q�8����!S���3$��	�g?�(I��I��4Ύ��e�Z���4!O�L�痆e:���dIW7�]-�t=Ӂ�|��Zx�D&�D�<�RB�*�\�����i��vY�����#�^��~��U=�Z��nZ����5��+����q���|K��@�/��jj��ZY�nn_��>F_��j1�a2�D-4�8�^�C����}�}�;]����+�����=�V��M��%�+s}�)�a����>�D�]�>�8|�|Hl��{W�D8xJ�ڇ�u뽛��.}���j__�`��j����U�\ �����Reb��BM������_V6��A<�Ň�,A�#::��9�}�*~^[[[���9,!!!�����b$2٤�%�b*c�VI�T�6�����H��^2��ԣ��צ������a��O�B���j�-�y�����V�r9wYҺ�O�oxYzyo��W�;>�566fbH+�szy{c
Y��q�(W�
��Gמ={����5��q͟�tM�uμ��G�u��t�\"�kl
�_�����<�c.���:J4�~)����ԝ�%g�Ui��2V�0^�]��]��uݹrk)޴�kkkT��5�ϲ�cc4t$��){�KJJ����2���R̓'��o���dKƜ���s� S��/�~F�<�X���2\niĪ5u�.I$f���� 2@&ap�YOo�4E<��f�h�C������˛��z5U54D�F���cc�!!!a"����ٛv�F0|G�o�kjlK%(��?�
:��~ڠ�@%�����7��j�~�M&{���I�P�Io2��zـ-���Mw1hx�~���E��C[?q���`��E������{���V�Nm4��Ue��_TU
\/�2�y�gS6❥�[qԻit<'*W%�t<�:PϏ�\�;�_p>|��?2-.�zȵ���-̜N��������\�+K"�)�X��ҡ��'����sK�xvCLK5�{΅:66�q@1�9b���6��X��F���'Oz��s2W,�VWWw��O�D
�p.������^U뫲��4�����J�Weee�!p� F��Qe�f�,�ׯء_�0C���Ϟ��֖���A��)G���lM9�6��צ��VC�r%_�31���܊h¨� ��V�2��aT�)�����֝]K��ͦ��v�i���N�����[&�6":G�.R�A���\�ĕ���'��&y~_8�</�������>bn~$���S��1����iKJJu0b�����d��X�b�x��p��7�����ڠv? 9�bG�����4�l������2���.u��������݉9>!���3�<���5���{�CS���`����\��ddlV���X��'FGG��6�t��FFF=Ho��^^^�[� ��ћ���i�g�V�u�]]1�9�u[o�J�߿k30���h�2�%uN�T|4�_w9�J7�g���=�~�׼�'�j��v��l�ܘ�iUo��'G���*����W�,Vr1>ǟS��VI��E�Q(<�8����X_秤�=-���e��z÷d9�%�8/AuttT����雘`�(�1����IZU[���	��s�<;��E)��Df��Im]]��%��GI��*��g�����sB�O��I)o��Ӣ�ʬر_'���TcjK�||fM��E���������*��\Ĥ� �`*����!;׺��~�Dz�q���jsPHh��rR���}/G�ރ���Y�q��4��wc>n?�i�[��g��]��vb��Z�f�Zw����Cg�\�oF�${`���,�n��]߬U�b9��SX5���s�e��FCQ_�ǫ��}G(�5��L���O�
f�:���>v7�5��p�C1S�>�B�>���i���������g�	���_�\sg&s9v�il�;p�5MŃ�>�Q7cSn����^t�NuokĄ� X������Ҋ���b����0�?�� $��Q(|YYy0�s�#˒loo3�����L���Q �}����b;eā<�^�7d�(��&��Y1�U�����X�X}S.f_�zb����X+��/0`���Z���".x_��8��0x���Z�$(.�yǗ���ۙ�\'I�T�-��ֹ̼��{�s��`ƌ�{�i��A�S�.o����<� M�?���� �VT����Kwj+�� F+���S8�%]m�`��V�����b"z~3|�~Yw���S�0!?W?�S��`�fSm���!���(#��߿����:2��f�o�� m��Z�vK��[�p5ϐ|�����n&�tU�l��mZ���W���n�c8��N���w.֟�%,d��ɞ��	e�O��:��Z�z�=�P��Km�%�`����_^0�~`�����z���j^{�V�>krg"]0�g��W;>t ��©���B-�@��;����%6������%�j?� ļ���DZ�s�|�B�!g�#)��ѿ*�s.>���]��􍍿}�2-����XD<Y�c���a��e��ʬoT��G��6�]��ր�Α֭㘰�lj��b'L�:#��Ss�F�Cf&�Љ�`�W�ܾS&wb6�`��o����3zY@� 4���JbeNTfJW�A��nN6z����{�3���������ס�[82k���w�O8����l��Xپ����a;vG�\KG�r^�,�݋��K�������Ӊ�N)��O�ą9�+�n�U��� 9�}{Ǡ1� �c8bB�^�y�������9<�M�ʚ�WS&�-w(��!�C��_���w/������׭��d��dG�kCC��W\��sA�����b�`=�^/~��93\Қ����G"uM��J��6 w�	�� �>�d��b�^1�#����T}���dۓzv����1}�ǆ�9DU�Y �J�F�@�����g�z������s{}�yF��}�e]��s�{�NR�r�nCg�9Tt���e7�%-��$��w��1�����G�����o�%,IDz[�K�l�����sռ�+�s$~�y�mۼ��ڑJ((�����.�P��J�4��@��A�����צ���5�x�L��}�+��_>���Ko�!�*H�x�^��&��tK(AJ�C=L�z�3�o�jP=55���[fG���Bv�B�~���E��'�@���2&W.)����b�ÿB�!U�u �j��m�p��`����x̻%�	���{�-^���j��N�� �v�"���C���Da
*ǰl��ܶE��U�Nz^ �8��b�:ēp�J(�ʽ)���6H��Kd流^�qF{z��x�yU:5(�Op��l��yG�epVG�,\r�������\˴��\3����Y�����XXw�M=NZF��ax�L??�Yx"'}��.hd���ٙax�9�}�6�:D�q��j�/Oݾ:n��X����pFoȸP���K{�����"�ןB)���J�����߁?J>�eY���|Ja��->5���SH�լ�3��TLcN`Jŧ՘�*h�}��,����uh�fS���cJ8*��
��,b}j��S1�ו��@�f�!OQ��t$�N��(�i##���o�W|z�G�w/~�]Y[+`����~RYYFa�p�CM9�2�+)�
��f}j��高�4�3Z>�|�۷;/�}����nN��GG�/=�ɕ�p�tn�0D�P��MƼb�}������O�1ۏo��9v�#��n>f!���f�NA(Pg��D}T���5"(% ]��tw#)�C�t�Н�����
�����C�������,w�=g���{ν?΅� �Qѩ�y���%��.ؗu����l:سF5W@n��Q!-�tp���v�����Ȃ�M,F-�_.�\;��2�@a�\U�S���g� ��7�wD���AL`o����ܓ:tJ�DӾ("k��n��7\� �ˬh%X,�ڼZ�}2�@�5㋢�L0��ds��t��aW$M�z��j+�X��擰!Wn��|�6��I6m�G1O���N��[���K�T�P~֔�].����Sn_v�E�I����7��8Q��oul�\�X��v�q����
[�|!������Kk3�(˧^���^
�5v"_�^�&:���n`[ٯ��s7ZtL��V�V�vu�����VejE�;Et���n�D�*��E�~:gS.�*�vn;�d݈�������y~��a^4ð5��6��H������n��/`FJ���������Ɩv��L��:��!����<�`�vg2�ـo-7�Zl2�x�cI�\�vG��=�f_�w���0�^���C�:!��k�̧�ygS�	#Ī<Gq��qT�a;��'��`�<L�FD'f� �S�_�K�vF|���[�<�aK�����nU�$�m����G��e�V4��A�ʙ
�#�����8��C^��;�p}�L�xmI�ڲ��Σ ��Oj���/����u_�t�̯���^3t "X)p���h�댑��Z&FFm<ȷ�!�o�Jѳ{QWXB\��:��#�V#����)��������}/&cHX������s�4���w1w����vW+N9K��ۚx��^kb{�������;�t�sw�+ѕ!�5^L��!T�d\�.��.���w�nd�r��y;P������=�-�^��ր3ـ��'5�A�Vk�^���h��Bƭ�Ϣ=/@M&M�I��q	�,3h�F������I�ˣ�ăfl�y�ނ�3fzA�������E�XJUN�C>��?`b��%��"��gÕN��G��l�9�=�gr&����O�y�[��������\����;j���������w$p�s)���� ��u��W�?��kW3V�lV�w��o�`;b�[��Z�k���Պ�|:��&�w��Ua�n8z4<�(�Θ{K����7�]'�+�2�K[̣"Y�)#���شj�*����GMG��.}��sjն0gq�9Zby�0.����4`���^zO:'R�!-��Yɝ��鄟�8�H�׿K]��	1����������;�� U;�9�|M�=��r_#|a����@�8�?�<��W�˽Y S���cE���Xmb_ns �Gs��*�̰�VR��|�Km��zl9��	Z�|Iy�햶�QqE���z�
�e�r.k�U�o�2�5��"�sӏu�g�Xf�}:uA�3��5�Q�r��x�����j3s:��Ȋ:��K�a���ނ"XQPZ&8^k0���z�� �a�m�<o&40�mx�����y��̿$�8��S˻o: 
��D	�ߦ�Ol�����������1�5t��۹db�!x��Ӱ�$�I#�1ڼ�V��3�f��}E<1����턋E�d�1�.�j!GY�	�43�����<d��q�H:����6IE�>�h}{1�}}��b�$_�" ̺�!��u�|� /"���3@�b��w�hq�:i���v�ECz�a�u]v�B8(�u�7��e��zQq�.k |z��Ľ{��<�Zĝ݉E6$*�s�c̐�}��D�2_1�P�m'/�#����?A�+H����B<i�0p���d��a��,�D��+�7wT�|oBz�>i��z��[=�<����|(��F�a��ۈ2�W�ͻDlY����{/H�@<�r�tS��E�
�Q1-B�BE�`���^���ܨ���o ՗7��j[tX1̷uTE隠w�pr*��E�z�<��3K����ET���Z��t�?N�˔���yM�u�`/ix���k�C޺rB�ϊ�	t<����	�HOn�%�֚����g���x��D��c�59A-0��`0-���[j��\z��r9*oF�4��/}�"��Y&9~o�8�>r��PIs�ǟ��������ډ"�X�)�!I���f�~�`����ǊP���y�'����A&و "_aҒD=�e��Vhm�D�÷�W5��$H1�7Rd6:׌�o�sl�Ti9׶���Vo�]c�k���Hw򠭼�@���(nYF0�(��,����%U1ES����~���7�`T���N,�<?��M��:�����N�J7Ӵ�86�Hf�\F��v��W�p���AB06����`���C�"��lH�i�켩����4� 6ݼ��p:�ϲ�V�xx�Dz!�X"��cK��L�,���:|6RTO`VC���$!I��ZE5��N��̾XɘqsF��;��;^P�����l{� ����=����4��%n��Q�=�Ţ���5C����m�(�K���P�U�{	w�3�˙8d�]�t�E�e��9&�i���.�mɷ�P"��l� �Pn���35�q�7A;�X���e{������Ļ�`X�C�a�u݈P��K�l����7�3iH�!�)�R�獲4���0S0���kΝ%P�D�4ܝ�q��4f����HP`8`��8�q�r+�BTOZ�%��_Z�c*��� s:���w���'�V_ ��kp$*��=�?�H\��@4nvb�}1�����%v�h�$�A7Kb���|���֩�&|y�F��b߃�ȉ3�Ka[Wa�'Y�^J0��ޏ�|��@o�='����F�m ���'�i�lh���m����Ⱦ���t{�r'ه���S���K��)�7���g�i��|<s`'�ksߤ���m���[�Xe�Oi�woK+�]6܁���,=_�v���Ж�a� �/No?מ�@��˴�7k�!�v=}�c�rM.�B�[���_朲�)�48�4��=�Vg�r�P�F� �Ix��,k��V�1@+** �9oO u#abb��3�nѐ/���)��������FM�w�<��l���"�\�$7��/W:%<q`CQ�h||���3�6�1��L���G�p�	��,�ӣ��8����2`m�����+[M��sgff��ё�F����93�Fo�_�Th�����G�	Z����O嶍nM���P_�>���GLFX2WR.��0���bگ�(Z(����Rs�Dw1��G��� C]��wC-���lɘ�}6��v0��e 7M5�w���īW�Jp�,��+5��\M��+�S.��5��{5�BDo�Q7�
�t�TJA=h&T��L�����5N�T⠹q�lDC�׷�,&M��7N)�Q�[��R�&�,���j!T��G���tp�|�
��׵eR��5�H��!%T�U�fĶ��8�3��xh�	�]�@�%���*�9��n�le:�`������}+�aNs]���;�**��c��8MY=������5���M߾)^�"=SRR�����ʉ`t�n�I�<��S���X�[��ߨ��e��{ye�H��^G�G�+��~C[��2�ك�o��i'�ⷽ�Qô=rs?�^.�aAo�7Or�[a�^����Z��Iه{��|`h���f��3��So�}4d
���4�srr��(�9�'�ΆKQ�����k�//�� �aJJJ�$?S�xDMMM2����P��|Hn.93���GZ�O_��w48��;Ԡ!]Nb�I���2VVt���V(�a#=3�%.�f����e
�TTTҳ��l��i'��]��_�BW�u0�������û�X�e�;�y�R8�~F��A�c�y�K��������3R�{4�~��I�:r2l�R� PW�cL�;T�]/�&��&5E׍(�&!N�{��~������A�/5����{�U�#	�#�0��Y��z]z��?�`R

B�~���e��fӣ��uG��O�s-&Cd ��� �����.��;8��u��B(�TW������&t����-��(�h~G��%��}*��2�ŝ�خ�W�j��7f%X�{GF0��c�� ������v��ܿ4��FYlv��'Q�x^�����\*����:���*�CDB�����������*\��<�?o�ב8�f��F�[�w&Ò+�=�yZ/U,{��?���	Jz��������������â޿C��3���L2p&��4h����x�&���Hk�(z4`���l�-]]��[f=�	666���.{�@T]�?O0[���PQ�J�+�X#��9&M���fzO#�����]��E�Ǟ���p!�Z�E�G�KLLe�&�f������	���ա�� (w0��9���x�KB�&��r�"��WG� �[,Ti1y-EuuuE���3H
o�Q��l�/<�(�f��颅�&�ѻ�,��
����1[�V��c��[���AH:�&���/h�l�x~�̊�^�ˀ`����i3����̋�B�������y�-읜I��Ybbn�t��F��%����@DDTf�t&��\
|��5afeM�4S�J�o"e��c�{���R�k{xx?0�x^�"���ёU��++���SC��i�f�p���ے-V�T*#@C���U�B����8��67+��� �l���͆q"��E�)��/8^��3����2!�
�?9S��h��bp�	�G=(h�]��������R�` �*sY�|����	z��[x��Q;<�i6�
�\X"�C�`fo�5����ТPW~P��ڸL���R��註��(��L4�&��_�PNO�4��ޙ�C��V]�i-�>��F�Mg!a�}�U o꾯U�S��¢��VcC���/>Z!$�?a�
�>&�{�i������R��O�U�z	q��.��/=˧Cs�G�t�`���x7�������K-q G#�I��ǈ
�&\I�rU:��tʪ)��Ddd4�?�V��G�?�c�C{���@�h#��X)W���z�YO�_��ڎk>�y�X����D�tUPݼ��6W�	�y�P��aAɤ�ǟQ�RO2


�`5O���zaJ��/�������پ��u��·Sk)G��ϨU��.��*��[�⍬8�v��[�9���3���5n=��+1lV��N���Ȝ'�S�o;b-��#0vt�aptb���|76�‖��
�|��7bʣ.��!�����a��/>�;�#i�������g�C���͇�X4/	��}���g�����?jV5J
�}yq���3>�+R��C�ծ�L0W_7~��ZFqlB�׏��I	%wo A�aM�s1(*+�>8�oA6��i*��.<��'�4C����I�j��Bb!��{��O"/�h^�k�&���$����(k��]��}��P��{������/�3�=�|}7}��R�sEzޤMu�㔌�$^���� ���r��� 㓷��E��R����@�����������NWz
�wt��h���#"����Q�OW�����絻m������B-��9y�庭�`(�����`YSGj <4�/}&ff��+1��&�����_�˝m�{��ũ5%���J�2=���%�'��{�2�� g�)�QB��"\��X�zu��{��w�qn��Z�8m�̡w%��Ws�>����� ߻O���|5�Fm{y���n?Qoq����������[;^��ʗ2ɔ;�c����/�2�����6��u�L����T��TiE*�F���V�}�%�\�1��g�]�r����s{ŬH��t9j'z��jS�Me����r��(!A��τ�Oz�i4�200߈�^]y\\\|n y7�=2:
'54}�?�.���.�B�?67i���H��g��>�uV�\�T9���PR�Ύi�Cr���L\��"T)������C˯��j�O���'Ouxt�â�[�`0;{��xU�㸁������q�ͼZ�xh�#cc��lf>9�π�H���DB����p���-�6d����
�=������U��boR��N�x=>N}�I��k�9��v��F*d�����M����O_t�Nv����V-~Ҽ��|~���U���m'V�⋙]�N�^z�y#�dO؅�����pl�m�	��4�䱂#��%<\
p����ϙ���!1��o;�S���<KsZS�����dnp���<�u��� _��'�6Ljjj���&�(���[�ᓲ1��<<�E �ew��1��&;j`����=�oT�l�������x��Lƀ�PO_���Ux�0�g��� �� 8���%�c�W���:::_L�V���S�	<K�܏�ɜ��V�Bj$��u~��뙷� ��%��:���KћL�8!1��X �#�<(<�y�Ux���Kџ-ɪB���Eک|"̪��	M#��Q���Qx��A:� O�<%-t�]r!;��v!?�-�|[�3!�;�RT(a���ܚ�҈��~�)�X}}�z��̙��B�~�.���������D>v�{��qS�06J"��$0-D�Ĕ�~\��� @�\�uEWf��}��/d0uc���C]��y�����/Be�*0�#��;��(D���Ôxh���s�&(��{jJR0����'5�zcC}�����V%~�;�����Y���$�*��i��.ޝF�<��HIL����
U*���6��\5��oFw�f�0�4i���E��gYq���G���4�y�fI�����!��\_I���1����'3�އmOʻ��veA�+<4��+�$�3��n�R���ZE��U/�MH�5���h0���Y�=i�%[�9u���46r���~����4�����,�����3�|r���s
��/��!'ӈc#�c��I��I�扊��ʕ�j
?���7 >c�+��g�g�O ��Yr���9\�Zg^��39��!�L��Ԕ�F����]-�6���b�M%����*��~50�#)�ƩS)R��%�S�~�������F�b�B i�̬9��yޞ @^�Z�w��u�J����ٙѤW/+���7�]MM|���ʋ��^����b��6WfE�fG�pe �IjҋR���H��>K��̴gӻ�M7�}�����Z�D:b}���=Pn�Tݜ�v��`Ѹ\�k%���=S����ՠc�1/�Z�w�@�Kȸe�&�xm����6���mt{t/>��k��̟�0A�����y}�\����!U���R;
  ww_5熏WrJS�q2���Zp����T�ٙ�z���p���^�LW!kW��q6F��1�(����Y#�����TK:�ˀ$�o�/���I�5��r6m������.c����b�v�"��~��O�oR� �#tւ�Eߗ���`#1��	��%�j����+;�s >���m�`wr��Z��$qS���5
��.��,C�y�f����XQ�9*��k3��|�=h��1J\:*���t��4��-0rd�e�2;c��d��+�@s��F�>�_���Q��Z��kʩx'��ylf)'.��S����z:3ͳ�z�d� �t%�i�{ՓS��(�FM�x���	����gG��I����3�H"���qME�%C���u�тg�o�j#�HJ�̮��C�z��5��\Ey9�泋���8�VkS݂޶^��8Q)��杢�(���ė�Y.��8�[Q͛��9*^����b���K�����Ez�ؒ�F���0O���ic���Ù�G�[M�{���S��nR(�-���2�x�V�z]����+���ܒŚ�H��V�]�6o�������w1���oϳ>d��W�<KՈ7Dzt�{?HL��@b�~�̀��	�{��̸.�����6�*�qK$,��zT�4�?����D���L����e~��X>Ρ��)���ݽٷ~2p�I�<�2�Z;�N���Ѽ.�x>AA�~�~�"�]��b1� ��V`dN�HpOyJ	�~~k5Ɖ�q4�N�턧�P�Ÿ�T�(��3TFv0�.��3LYH�f�/�8�|LH�5;�l$�<�5e6�B��a9>�p|��l+�uTO�l?N��o�n_��+�1�~c-��bE�e�xrc�
I����И���I��ٌxқژ�4n<��=nXoW�՝�y�Yuc��?d_B~��Ljt���j�V�թZ�]�H�s�+]��9�B4�m4�g���I�_m�DT�%�=D�<qS,���"���o\:��^�NRR�[�ưP�߱����QQ���o�i�.Q,�U�u�{�<��P�?��D!yi��ug��d�ր�d�u�dH�*�qT��2�z��l�Q#����?��ZS����A|Z���<�,>�剚��*�]{�wUH�R��!z��'4��?��WȶπG�0���D1^���˿����0e�:و��%�����@c�镨�M�Ä�Y�G]f�2�iXZ��S[*�u���[ݸ,p���ֆe�������c:4�;~�ʞ��'GFSzy�5L�Z��I��ƒ�%���A%7&���^t2F~���;��r�z�~ǆu��ܟ��ntB`�oDw�3���=��.tCk_��a�2d���Qϧ��J6�!�k!�|�hɽf���4k1�˙L��p�R�Kz� `��rވ���N�Шs>�د7�X��k��kWB�/$�,�`�Ef6�/�E�eK�X��BC)���$����U	w�:�������w�N,�����j�n�ٵ~"�|���x�e��B��+6����
l�z�%���1�Z��N�T�$$����t��Ͽ~�zj���5Q��з��m��Kz��ބ���:V��cB�x�B3�ى�ڔ����o]G�u5�����R���Z�E*��+AB��~Y����ݤ��Y���,���8GՊP�x<�("9!Ƶ�D兕��@ٓ�D������C� ߾o��IW��>7�urFo������_��L��Phml��۳JNH�-���ĨYf�;�r����O�E�5}�e�����M8��[��WT]%N�+��:��eѦ��p�Kv��ܪ������m��,�-�] ���Ҿ��g8}"���"������E��y����-�%K�6�$�wv#<#�%�s�߄�2���x{��˺k��K���N,��<(0��L(�s��/%��׎��n��#PD��	K�\��Ʒ�LQ���7�%a~�a�rF�:յ��ya>�?~Ѥ�-�HO�ˢ�g�k�O�v�/.s����}vʮ����\���m2��r��&)�*���K�`�xm��Φ��㺅���
����=ŋ��=����U�4��`A�*�q�����������D̏$����*q����
��hc�J
r�n�V�6�x:�=f��h��-�:"EI����ol=٠�oźk�XoHScmL�g��(�ݠ̻c�*+����Ήz?���.�?���j�Y��0|���k����O�yZ/�Iz[�Mg��Y-�(�`\2�'�@��e��jb���;�3�UV^_�Ĵ;��U9�&�W*�e�:ː��b˃1������v���C'
�{�$}RHZ�����x�~�[����
^aB�8:~����)����(��VUQ�'aگA̚"̑�D҇9�����!L�Cه��d#��zMvەcN�%^T�
X�]B7���.8�p�]�2���Ȗtj��(�(K��v�6�8w{�<Z��]_��2)t69w<3��{ߢl�w��ۛA���yr��rҽ��DӚ�0�����]\��ێ&I64ce���	*'�Z�T�5�̒G�*�o%J����ok��<�r��%�	��p��K�.�Q%�7	Tu�d֬�ov�9%�0�d0]�u�7���� ��U�/�.~��
���]��`F�������� ��k��Ke���D=v��S�*��
�m��hul�-��hb�b���G�)I4/30T�#.�>����؊�^�q��� S4�"n�~���Tg�b?�
#�]�J�/���q˵�ڱ�'"C?��p�ג�����/;�c��qE\��v�%Ú�#F�y6�6��s�
Δ"�����S)ha^Ҍ��5\IE�99��(��}S|}/��O��򐈕3.)��Ք.Yim�4�BI���W�ꤸ	U����<�	��y�#1��*���Vt��m���"鷟&;��.J9{�!�O��j�f$9������^S��E/0����a�]C#�+^I%�~2���^0�h��J|
UTT ū&����efM�HM�(���i����6o�5�$�o�Yq��F����{yYI�S�:jj
�Y���v0�����U0��v�̨�ӂ�0���$5���d�5�α�Z])�-;���o�9NI9���#x��3��87��ܽ� 07<�`��D�0	�C!�e�˜@s���������ƵЎ��P_W��5Z2��Ӛe$���k�މ�1��k��g/7շC%��@��4��e�����J����p�!+��4��+j���tوh�(��+��Sq��.J�?k���*/��/',�޶tswOV�͒f&��Ǔ�J�r��/}~T���-h~`L�%��8v��F��!k�eb��,N�L!JD������c鑆]IF�^�:����ک�Њq�� N���wƞ/j]��r����aYE��ܤ�' Q����^Z�hY4�����uUU�g2w@�N@�G~P���Q-!fDa��"tU _��ok\��[@ ����B�e6fԒ���zyݧ��ʺ�k�xaw,(;����%���AI'������a ��g�[n��G�v8`�0c�ߢ�O������OM&M�Y��z�B�}���$�i+fҠKk�@�3%�%P���[JOot�!}��4J]�Ť��?��m�qs���ʪ��f���ZII�ڶ�j+��� ������<j�s���W�p��7���/j�����P;�o��0�e&(l�J���vp�����D�V|Фj�x��+�[mS,N�Ȁ��=8�md�G��G��o�}�Jt뇯=���?���3_5r53*
�Հ���@ZZZوzVq��7���u�t�����t������P'�������1�<(@hn��'����2C���L���Y
S�,w��S���$�a���ϋ�����n'���Y�1�G�HhB��ˑ��@�I$�5�w��Qp�	"��5[�־0l�cVFrD���^�S�lJ2i�L�!++Fd�^��o�b ���|��?0P~x���9,4�ն�u�S�X;:�����q� ��t�|�"W���f�I��[�[N��9�+n���D%��613��%VAiiĂRviI	v� ��-�^�dd&@ovX�����6�~8��#��$���jr�������ܯ�����ͽ;�[�[��>ًipxw{a`bj�ˌK��,��2f�A�`�TO��/ǿ���c�P��w1/ L�%�1��F���y�W���y�m��D ��.q(��(��H����t<�QV���7�P�p���)��yv�U]��B'7qT�/��/��X���uz����Hn���A�Tk�<<�!U���5ۏ[�}?�==�RS�bbb>geQ�^�7.�*�×C+�f|�Ԥ��	�����<� ��S�Jё�!ߍ�Z5�U����	��')�:��D]ǵl���L�l^O�A�[ʝjv�������Ύk�z&3;[�]���K�^�ճ�i���O�����ߍ�Dj��]�{z'%`LT��/����v��k;}���1\rs�$c�0�@����f�O��&��i�BJB�����fY_�(m�����+�4�7�m��0ah�W����@����Ȉj�o��z"�ʈ�&$�w�� 7��(������1�8�HR.�����,���ϧ�[hA�LIHxC�� EE��x��o=cڢqx�-��i=ф<l}�F�Fb�ԙ��O�' ��b�4r�����R�2Y!�3ŎP���O%���K������f�9�g1"�D��x����]!n��m��-]�Ny�w������Yb�ya�G߹����gx�A��W�0I�ߍ΍�/G��g�a��7Zeh�j�w�=�ᙡz���?P�(�"($���!�����m
�˦�rJF{����W�]�I ^1p�bM�����[n�@����v�Ғ)2���=(2�3����"���������&�O��ub�"�t���X
��Hm��N_�T��$Y$��|��$aπK]x��_��]���x�J�oB� �iw�s8
}��f��3*�����ʹ���^1s"�V�X��c���-O.Q7Ÿ��ۄ�W�s��}������6J�mN�<�ɔ�%����w�y�d,��=3\ �(�����ڢ7�Q'~c�z:�y1�j=��
t����cL9�Hoo��~Π9��Ą��ef�/���%eSۇ�{�?9yy�f{���d�k�I��{.]�_��^+��D|v��
=�h���p� ���>Hs
Fп^-?F#7�ЅEx0c�||�O2@&���hw ɑ�a�Չ��\&��8Z�M����p,WjWQT467/��
H�����Ͷ��!0������A��c9|Y�R�4�2���Щ�ˈm�����p��i���S��E�U���ۄx@w8�I��'?na%u���
Z��}�<L��T��b��<w[V���ܔ�Ƕ�588<[=��r؉Oq��ŭ�N��;���L�����[o_�/.и�h÷
_jKiGB9i����	�A���%6>~�eB=*-� H�nD���0��ws�###�^^�E燇��K�Q͹~Xn�/�@f5����sA��߯X���!(�PB2̃?���	;���ɬp��N~Q'|�`S�����z{ē	!D�?�A��zg�\�X޶']���jӳP��7��IVƤw�]	�;}�ޖ&d
����˛�^Rl�g{OAZb����M���[��K�� �2�6�	�&YteCT��O�a�j��t~@	C��67-Yq�ӈ,�N�9�n�D��2�ﴵ�������� <!uf��^�	�%#��y�k��f��{~�j�UzcSSD �����T�&�~���AQ�lҨ�d`�钇�;e��Z��r�:��5�������=_�vk�����v�{�z�ᴊ
c;���^^���C���!?( ����81;��%����x�g�DD.��Vڋ�,�89�)��*ٱ��������7�kqf�\ZZ�=�+�%���+��M��(��s�������Yl���l�Hrq��r���G�1Sa!v�mT��}�~�e�i�X��go1U��M�C�G���茄�ͤ�zK��D�H҆ho]x��5ѷ7�in����LJB�ݙ�n�0�ZH��gh�:�3NX���Ddm̈́7� �TPP���Y=~���!����76Z6fD��Evycc��~�%7O~gg��E@I�c����2�c���k2�H�t��~�jHH�C5��i��������m�- �W�#�y��?��&S9&N����0u�w��K]�t��DD�����D���s�i���S%�c'����wq��x��Cfuu��z��!%��� �#��WMZ��,M�`���[�B�`��DW����^6!o'Y��Q#�o�w	�OV��ς�ȴ���o lXn�a�o�ΫT{>�Tg~���aUn�V�:��;o1Hv;h$���>�\�ϓ�I?+�
�o-�I_��Y��U�FnFg���`��z�5<���`J@Yp�z�-`OoS�3j�����t���x��3�b�t�cd��N�َK�q�<��u�SJ-�f_��I�@"(�D;��^�ᚷ�usWk*����%��z]A?q��ʊCH��U �R�C1�����Tj��U]]q@�	���c��֥���`���Q��G��r�R�E@���g�űlܯ�mtL>��P.�+��Dm��e��{�o��KWTPa �^߀�}t�C��9gF�q���r��˂ⰱl�� �ff��"��h������7��'�[H�9�K�
u�,E�|���|Y����QȪ�G�.b"�jz�?�k�/Z���Ă�Ï���u��觡�Ŗ�0�M�#|AQ"��`��[Wr8R˒��U�x"��/���m������>��8iw]����W���1|~�橭d�H� �X�oڢ�qJk�O�̀V:���'()<�x�4w�Xȳ(�r�,R��"g�gv;���Nͫ��4E@�@��W�(W�ӣ5�p"���/}ʗ���'�_m|����'�X�����t�i�،��L<�
p>jPO; G T�3v�Oxt���x}��^V�XMA���,دOP�D�"��y
c��Ky��)��+����bmw<BF�$��7�ݏPU��v��kB�g�/�$?�����ԉ� ýyG��`Եi����M9�F<�Br�Y��-���]��zD�ZC���h�GG'%���/�%e�))U�ү�J����옚*x�w���Q�����?uf�7aT�\�E�l�v���F�xCeoeDm�E��N�F9	8iT�&�ʒ���<�<�1�#���Nl4Ɠ��y5��_	d�$��%ټe*�:����,�ܚ��g�S�ǈ2+�b�Ŀ��]XRs:^.B-�e٨�~2
FKfY)<b�W�	rr.Z:�h�n�OB;���l�=~�b�Q���ᕨ⣷�o�L���K�����=Ou��i�'�(���?O �07�W����R���j>�vb��T��������̸��Bw�]�-@�ә�䰑 ��T��L�W�����:GM�i�O��(�	�*ń�7-o�&b�i�� �U�K?lٙ��1���/<�pЕ�u�j��e �I��b�|���لׇp�_�u�_��R
�XX2�?ճ+�!߱���cF�����ff9�?=�|���nF�1�r���j�	���R��0�#ҷߤոy֌��L�%g�F���Uui���z��w��P�d�B{�8�LϤg�m��Hf95Ӡz�q��H�%��>���rG]�e?+�Y�I<hc�V�o�珛L&J~;O�*^~�+[��kRn�[�D�;;��� ���[(�gj��:��� \����Ļ挀1x���?��k���~8���:���b?Q��?[��o��f�_�7y��G+6�$��h��VZRK��Ĵ��y`��nM7~����Mc��܋RU��mbҶ5����D�Cqw{�S����B���f�Nq��1C��������G�7|EN��K�K��Ͼ���&�ӿ�C�C���x���qK��܎�uӃ��d�ID�_Ơ eb+ܸI��L��Ebfa����EGK��%
qZ�wS���7��E'�
`��o>#Ox�$�s��0�w��5-kL��/��d�dR-S@�uI����L���� ^=o��I!��ޫZ��⦊*��՟g���n�n����ذ�]]�6���qO~H�.�+z���lߦO�+Ϲ��&��"p�q�j��O�]���$���	�=w�@��z��T�n���¶� ��lx�VJ1_���NE=��ݺm-�H�Lg/b���P���i��0�/o�)��$�'�kF�	b¢^a�X�7��[�4T�C=+�j6�'.���������Ί�@!m�8�צֺ���,ߎ�Vjן��xsA(���H>&��@J.�Z�l�Ӓ{��x�%�t�fLY��ES&2����=�֣G��<�7�xD�8����^���m��!_ڜ�ҁA�q������K�u�P�O硇��w�P�-��H���<�=�C�^�1�ha�P�=��W��੏ݓ݁3"K1r�����z.4�^{ Xo2O�iX�����[������ٽ.aw��6_w����!T��M �^`y��Y�~~�Iq�YK��*��pt��F.����@��Oz�rI���2g�^���58���ۻ�t�o��qV��bh2�-�U�e�|�k����w�v��Hl'���odw<a�m�YO�6F��D>��T�N>D�b5x���ѯ� f���g��ͤ	�t"�W��o���R�,`�&FU���e�ߒ�j2����>��Zu�ٯ�mBھ��l�l(���L/]�2��ʻ���c�4�e�9���t�D3k^����°s�;��M{O��a!��¹���D��}�?�Ly�6��e�P�����H`4]7o����$�+��`\�R5c�-���KOI�����z_�sp���ı?��+����@�t&U�ŗ���\3#-�<Ŭ5���f4C��Zwj��_pK�Jx�9=�D�&���-���>��"�;+!M�Wu��I���V����(�p�&5 " d�m��l}��|�8����z��r&��n��-��w"��	�=P�yx���;���Ƚ�X������Zoɛ���\W~X��ɠS��g�S�"	���*u�$4��j�	`q���7Ni�s�e��)}JPf�����Q�D��p��"�2ڔ%����*�ѣǟ�sz2hF���oߍ���IW��jm��v����̀z���%�̆�pR��Iet��
:�+��ݓr䃍���H<�!�.���D{*�J���%	�&����s�� ¶��t�����R5"RJ�8�{)o=��@���ͳ1W��W`c$���˾�KK˴�so�ʥ����=O�Jgmy "w���:|&S~��M�D���x���X��mr�4~����e<��5��t��"HK��vo�z�^�������jۯ��o�)-Ո8�Z񥃪�O�K��:�B3�?�a_U�M)HKJ�<�tIK#����CHKH�����t�42�4C�04�|��{��׵�p�>k����ޱV�>p�\1�n�S�
r]��H��J@� �?^��@H����~�'��TO�!��@OUS�?>�]���K_-�a�AfaMM�y�i�y�@�RB�U"����/'~��ק�$kTt������C	����`>B���9���)k��F�ha�s��D���.��c�`��6�8�?��7��d@m���\�"o_ך�K���-�z9rl��&z�ȅ�͆�x&1d��S'�~�$}.��]���LFlVק��N1hqd�G���=�P<m��Ͷ�SL��:��*Eބ�5�{���h.��[�(�n�3�sK<�S�5�����$%s��$G�-�������ڿ����>y{���f������2��S��vH��J"]�U%���
l�+)�����g;�F�A��Y�%�l�ɏ	������Zl�5j���ސA����9�%`�2l��
z!���?�F0^6��y�{�������Qu}+�l�� �.T�/�+0G^5F�������r���Ծs�5Ѝ&��p����eg��:ϥy�]E���s�h��o&�ω�i��>o3��"%��JzUX��T���=^���=�-�+�����i	\��S�(�|k������]��{�:0L���������r�0:6~?I��'[~��b�m��t+��%�n�[Ds��O�Y�4�l(zWG�/ך 蔐sr	���}�"G��~'����a"2٨�y-�G�D@����
�aE��ѩ�N�-,,]�����$ZT�9�����[��m�?��c%a����a9`����K�S"J�3&���	�jf�	-)a���5���ۨ7�W(!~�yF�ξ��ZL�w
��?b��ϝW��M[��	N�X�]8�Hu�T���N����W+x�JU#�"g>g�����;���A�bԤkb9�TNi�t?

�>�i�� 4n�뇝�=���E�1<٣�Dv6R�wZ�TB���=����)�����=��o�e)2��aI���[FT�m���be���tY�g����b�ݎZ��:O��b�x:�ޓ\�F�N,r�����E��?���(���5-��0����˵Hޡ�2�!Aa߶����k�0�k���1g��(���.�߰g��u���`L�\�,	�I6zrlv���M:��Z?��:W_%k���\\\d�&V��`�Z�g4��Z��_�\��v��	�X� !���3�p���626��o��b�8yx#�|�F��v���N�F�D@���(C�����(6��o�v���VM�m��q�M��N5��y�+�4��Pv}�Ejo����w��~mb'U���E�ŧ>U�]"�����:�����_�o�Q�]�p�P����=�n�e��$��i��4�WgNY����bTmAKˋ�����g�Y%ǲl�����2�A&ΔU���A���Ye��A��ಙD*�C�;5��������.h(b.��,z�<;��cBD5�992� B����1��v��O���$����V2-@�E^K�Qd���]��"��:	g�	�a݋����~�����y$�t�{���Shڝ7��~J���!W���8�@r��3�z����9Ogu���y�/u�������<��^$k�?^V	C�0��s�d��"e��B��8]�&��Q*�}#lX/	��^����j��ư�`��{Ȓ��7gW�;��.##�{,WT)�y%wD�	Y�F��y�yn�{�QP1C)��z��։"Y�1D����+S/���+~!���G�F��7��Q��Q}�5P���ڳܧ1� ./�;�H����]��h$`KEE�{�2�/��葵���B��<��MLp��T��1����4�b�I� ��V��,j�z��A�yX�=>�3��W��I�����{�qM�y��Ӥ(/�fq�tj���W_�E.�!�k��.��X��2��*���XtQ���Ʊ/��÷t�&���� 6�M�*._>�n��qE^(����a�fHk Z�i!~%��|0!yq~ۮ�T50 �ˎg�'OO�v�pٕ粒�9MZ�Q+	!~�c܇�uu����vY�K`f��ȅǙV��{��Pc����� [�uUM�\y�'��O>�/���h�bt-��|�(���TF(�8��.D
Ź	��~�`��D�ޚ �ڔ[1�`xQφ{�ʯ��PU�6�ǹ��~��]mB���㖜�2�ԃSSD3����������4A�kkk�����cdR��P�͛�ȎR���JG(�wT���_|s�� ����YkV�؁�Uacu6=��f�b�L�I��D�~��'��o�z�?����d�RB�Wy<ƥ��=�|1����~�3�� x��ᙈ0g �����ɫ�$̤�`�-���~�d̐��˭��M�O2id���� n��ｧ02��G�ܻ����&V3��6�|��@�3�
�����3@�oooKd�����������@�h��MV�$��l�����hH��͛7�L��-�/�ww��P{��4:���
���I*�J����u�\������w�`ys�1�>�B��Ξ���w�f�[���Z`�h�����/,
�yzy��\i�����fZz:�����Ņ_��A�,7�~�gBT�rssA��ϔ���q���߿*斔�Z���@��a|R�����l���"� ��,�C��ϙ#r���I��ݲ(KzxNB,�So�@��Ɏ������6_~�su_���um���w�H�ٽ���
��f���qs�������i�Ifz�jM���$i�����lK���: .U}�㈪EqE�/�)���8���ms��o��������?�����L,.��M����ALL�ŬUZZj֠?9%������A�c���Y5�^�)|��(�'�&%2��aV�����\��1�����W�)����AGGG$���k�`'''a�]�Ԕ��������9BU��&'5w%��wv������[Z(TUU�����v�X΂�)��@�3���q�x_���k"�qn[Ƀ'��*��Ȓ���Dq��ӿC�t�>{��*�g}bŏz����\�ٸ����bjj*��op�`���e�-O{,?s�NƮ�-�NL�w����)�ѣkb��L�;���(����,DFN��Jh�)���nE�Z��kF�b0\Rq��PU�����92�Tl����4Ry��������aqӂ������BM�G�Y��\~���-�Pn��gJ�<��Q���0�I b�tK�v���n�rgycЪ�ej�?��O�<�\���q�XP���]�	1C�n��Z���O%�I䄩�e:
D�p�����g��;f�W7G�U"G��V�����q�H�{��ޟ�vӫ�H+���� O�!kO�-��S\__+�	NĐE¥`����Qk⊊�f��W�g�v���C�Z���nnn��:��8����tt�~l��"�$Q5��o@V��`�@9��g���u�7��hC��&���vw٪�;�w�3�>a��:��ܔ�=����C����DC��n���.0��s�ow���N����QF��-9=�5�6�~��x�oj�_�K�������L���_�4J|;��;3�5A�5��?0��H��n�"v�a�d8�T�x�@��bUߊ�^A0����.2��X���ӈ��|��CS���7+�ȱ�Ԛ�tA�fЮ�&�}�1��**�c.�Dq1��2dllLw܏���k ����%/2�9�غ0r[;<OY̊��9j��Zm̨��j�ֱݚ ���)J���i��́W�)T�kno����%�y_�P�|���L�OPH(�Q�)�Q[[��~�I�����	O��6뀻�o��[%OG�v�/����	�A�>9����x��ݽUx��,K,�>e��ѐ��h�&�Խ�/f�m��|�%/��d�Y?��3�����GK�_������mb�"Ԏס������L�i=���Q�J�Bh!�+����M��٣�)Cܬ�X+�W�J��A����Z_o#8-�h������+2e��u���L={�[��]�z`m# (��솮��la�x�Q���qp���ZU
%�y�m1M�<P�L��yGs��S�.h�p�JЦ��: j�<�88���y��ƚ$�v?b�w�E/J�ˑ����G���I�B��,A���*jj�"��X�̴�
��/�4�]�(I�PI�ީx[�Di�w�b�{����(T$���@��Ƙ3���>Bƺ� ���x�Z3�����侢�;�U�Gd��H4�"���~���3�2�*�Ʀ��a
�[�Q�iY� À����M�&[�F�7�$i���RS��ֲ��Wa�ձX"�U�Դ�ܶ8�nII	����s�"� �#K��hE����-�z��m|'����a|K�bF���A"�sp���� 3�C ��A�$fUH���=�����8c������w��E"����g5�F,? �����2�2�J�e�`�؋�� �T��Y�"�m�i>_�>�~�h�|ޡp�0�&A���ץͥM��z��"%tG���dr�f؞n��wY��2��Y#�;���=�-��Uڵ��u���$"RE7�� j^��2�aJv�6��9Drp}����4J��'Ժ����
h<�H5��6�qk��u�5���A���G���	<@�-��cc�)��n�g[߿ǔ��J����2����w��>�3T(~�OK5\���`�GR����1�Y�����;k꫌�̗dT�L���IR"��?y�������C�.9(,�-�.�th��W��$��M�q�F���T��Y�Ka>Ґ}��8��]����������9=(,�� ���s��Ê�p_�lLl��8�3�%�1G�e��V��[�U��Kx���qH��7K^��<��V7�hY]X�f��&g�(�w�� g�b��刼�)�t�[ǁ���2$e�v!Eo��H@����e2�@ؿ��
v���ɑ�4,.�O} MƞIpҫ��k�������cк>��y��V�9�y�D1��7 ���}��i��2��;�cɹ
�k�.��c
Mp�e�RRR����j��)��e.<x����V��
VW!n;���+n��Xi��/�g�K�5��}��W{m٬P�R����5��?����S�?�ԓ�Җ)~��L��]��r�I�$�A�t��{�肾�YF��	w������LҐS��i��e�Շa+�X9f�<���w���꣎���ǧ�ܸ0i����!���7Aȣ3ƀb!� y)MJ�J�����ة�R�g�ǩgdg���Z�Y=t=_�s���d&����T>+/�T��F��΁��YE�)�<�Yx B�x���ù���-��Cx#���{�����f'1�4���G��̎F�OS��?S�u�{�2o�kT�b~�;ssh#���Vo�y�iP4��,C᧌�������%�5��9ø=�^P����4mS`*%�j�3��dY��T2�d��$rGb P�%r���u ��m@�e(�o��#�e4��E�KM�LJ_���5H�B��0^>q�����xP��#A�"B��뇏! ��B]�_�b����D�2�Κ`M׸��V7n���{�dZ��� JXK@[����j�O�z�1l�w��yg������@����ږ�(}�X���_�����o�&�po��|+q��?Z7Q3��d%i�����k++��=�K�� ��n�ܚ��"3����3�S5c�w�$�$Fks8ؑ�g���
��Wy�����Ԑ�޲^oX5.�At�Ï{���?>�-���@�Cj��8�+'�ȃ�[uqkϭO�6X�����0(B���sb�¾`�?������=�O���S�XN�Ǿ>1����Q�XqE�O�:�{������V^� kK���GkGT-����珟� �+�r ��U��e�*����j�+&�'K���}Y�o�0c�bX�
����n�l�988<s6v�� @���&�AV��c�adLz7�'Lʎ�i⧴�fA����
�bq!���e�I��x�w���FPp��N��Z�����r�{��r��w�k���6=�	�e���@���{� �J�~Rʈ�v�zn�n���kZU�'����R`��Ǔ��Bɐ3�j�6c��R���fϵ�0b�u��uu�� a3:I+��XtK�_���qu�
��'i��	R���`H}�+�����t맪qILC�Akڭ��DQӁ��|�P+��������!���m�q�a��f;8�)�.�`�����X���y�|u=��շZ��[�Sn��8����7"�P��[��S��{�I�*G���O�w��S�M���pd�i�v����s����#�}Ä���r'�����h�4�$�����L��湵V9c~I)����h㼖��߈:��<����a�pu���@)����y�\�tf?�H�HN�#��E��*��x�������c*������o}`�p�Ռ}Ö������ʯ��澪��5��� �A.�r��5��0uZv;���%l�yiÝ"�>缹oUJ�V��1a7p�#�!��/���������r�������8!��ÁX�6	��;*i9�S�Ï��+]�$I���S��=2Y��>U�c�|�����z���٭��b^C��n�TD����v����=��N�X^���D���K6��$E�j��&�t��JJE}/����i�̀~����Q5R^�Ԫ>8w��W�5��#���J
Y�[Q���\ݶ��eX=%��Nu�UO��*������+�-��`;�2�ZeSj��;S�����&�I�����@ ���}�)�"˚�ܨ�M"�L���.s7����z	� �;�ٿ��q���f��G;��q�O�;�ܳn~��J���hS�QH]w�A�9}�`�!(��^]��_��)%B�xL����FԿ�׭�)��A�Y����am7��B�/{��4Gh{[�-e��t#}��>�QjU.?\���ܭ�~��`�9#�;"�Δ��D31ęр7����Q9i�6�ѯk�$BL���up>����������ns:#�-@���� ���X���,⛯ީ����D��_���'�)��,��#�̀� ]e��c�Y ����Ǔ���I��@�������Td���`���I�z싛����J�`�~��2W�h���д����,�w����w`|���o&��&��+Q#�p^��_�Q���=8趕���Tg�M�����9Dt��a��S��ط`�������pR�j|<n��Ƈ�~Ԯ�^�y�c�ݾ8��$��N1�P��%vi9*uun��Z3��6��+�Á~yQЭ�+����E�v.W)~���)w����w����=�?KwA�uԻz2r�Ky}7*�#���\��/����ӯל-�\ 8�+�9�o�?U.�Z:��ԯJ��`�*׮Ы�o7�����>{+ q�j�68h�+��h�I��{���ǵu���#	�����b\�1J���c�]Rf�/d/IV%/�k$��F���"0�<?C��E��qI������L-�����!�<~zuC��3�����Զ�^��xǄע{0�lL����sU�����w<ԻM<m�`
[�%��쑉.�rU���#<Nk���ы-+��Y����#���C�n֛q��n�H: ]{��N��ꁸ|9[����j�u6ͦ� W4�W4�;����
�w�!��s1�������։5��!%$�5gz��Gp����*�Dg�LJ�Uc�Q:�+��Qū�`�k�,ܸǽ�&��;B��m�j<MU�>�����Yub�� ,�Qnl1�u���#p�5X�@ �?i���0[���{�g��� h��%�QP�7)_���٥34���E�}i�v�����}:�t=a��ieqɑD�Ȉ�����V�`j��g6�W{#pX$ ����h�I�^�5�X`��f��E^���a�����[ߨ{&�'���5eL)J�-�(�d���W�W���Hh�f��eLx]����L8�7at[�E�������Z�¯�k���T��(��kN<N�m����i�k����݃�%���7 P�������̴DK4�2o&��`R5<���2�i��d�P�@�?�-�e�-!�d� f���aLKKå�$�>����H�/B�>ڷD���Eb��q5�jY�V��-Bf'��
Y�[3yyjr;���pJ��-�Rk<q�'؅y�dh�-�����`���qA..��sG��E�MM��X<X]��mѴp�Vȏy���ڿz��3��*���?�
����&=�/Z�Y��0}̯��B���lSK?�L���
J����G#�߷NT��%�m!����E�8���d����Ak�Į3�OR[_oQF
Jf�	�|W����s5���n��.�^�"K�Jzw��vus�<�.���W�ű�u�x���ײ.�+9s	��Z�TF������#�.�~�W(	
����V�'tp[��©)Ю��p?=��
�݄��$c=cц™(%g85M�7|ij�6$��7d=+_0�$gL�B�.;7�jV�hp�%�Zg�\�0aE��8c����|s���]��0�b���c^�H$rB<%���@�ڎ'��'3=Zu}�cJh\���){��U1�{5 ܦC�lr���+��ȧ�M1;��rtuS�>�E3cO!�:�6�D#**
�_���5k|��ϡ�k	� ��->?j؍�X�TQc���z�?��/�)��"Wh��߿�����ˍ�G��{����%��Bz9�m�0�5&�=���! Ѷ,���2-�L��O��������Xu��mV��VD\��6�?am�>;��x�}C�,c��\������Q_�c��[����737G.D�>}I<h�"Î�����aȔiI�f�|̊�_Z�>�B��>9��Ļ��Vh�|�$��̚��U��-ѯnXprtv��#v�����s�%}q;�� ZFn��l�$���=��P@i�ֆ�s�g\t�-Y�O|��p�E)T�5���O͠]pʵ;���+Ӂ�����U��]'�����jXr������ۑRU9�e��(�=��հ���h��FGGw��Q�ϔ�����]
��!�#�@�\�mZ9��L}�N�q�k��ܜTُ;�浕S���������v%"�-��o�L�_�)/g$��<�n�k��*wIX���ذ:������{���t��Y�]����A]����j|mF�L��ONN\Ere2G���H�Lڒ�{g����qRQY�iM��Y�PFH3TVV�S���{�QCzV]��b{֎?�W����4�	[>�,��J}�{�fp,�11�߻�R�ՐeK�^���w?��t��\�����s�V�ߡ��P�u����{H��j"���/��	�?�@!R�|�:�
6��F(����p1��W#��J
4X�'�}|҇ʭ axXDDDA8-$��������.��U�[~��o �l΋��3u�;�3:
d���>?^N�s��"ejY�4X��h��D�}0����!F�4�y�ćW�6�K��Ȁ�A�b���K����>��9GAd�xkk��U��WanT#hf�7W���0u`�a�F��B������ �I?,�6��nv }7���W�4'����e��J�4Wg���{j���V+�MF�Z��:�[�+�����׏٬HL.(|��:ep�8)� ��} e��݆׵LP:��j��ݐ����5}+B�$� �8��kZp;�a��$�W���$�����K�!��3�PS��jV�{�m83� k�jKx>����<��1������E�,w��T���"*))���]@޶� �V�j�*���P�US�虸`0_뢳a�?)m����/a��.:�D���J���Eg:[w��W�7S\7ɫ��,�,�N�n>�	�N�qh�-�GH7O�Qz���;*�2l�u���`�v�<����]o�;p��};����'��Vw�}� ���G^�,&oNO�X��^$�J�Zׯ^��s��c�c�m1 ���<��/���z.�n,2v���qK�Jm�w���G]��	�&����H�ĲnX�|QH��/����X��0f�D>gzl�G���o��lx)�o�H������;��U��@Ā��U���\#�s��x^�� �jC�+�T@P��Hh�:6��Z��	���V�t���Ğv���u,���mr1��p�6'2:B��Hn�k
.�"�U~gE����+�Џ�P�4�W�*�K-_��lq��-"yA <}
,��1��݆�1~UQ}�Q7j���w�� �Y�G�Z�����"
��W�!2�TL�b��fڶ�W ��
�`G�En����]��>q���U+%�E��Wj�i~K��"UQ^�?�ʙ#9��#�0d�����F�~^V"?
�F1�K����}�#��M �B����(HDֺy��C�TlK���-8�O!�
�����Qld|��2�II��yq���/�o�����^���H�}�Aь�t�~�Hƴ��r	����w'�)���tB���Պ�_�T�no����� ^ �����w�[n"���S����z�hZ��Q��G��" ���0�
3z���
D���;:9�̎�B�	��2s�}�=]��g^�մ ^'�`ȹv�����8�F�����|��oҠL+<"y��IY^�?M`r��ǋ�E���#��hQN��mY���C�t��I[��!)��7��ů��Po��ǩ�����1 �n����;� �eQ��k@�c/<O���(�ZR��=�ވE�7$r$��u��i�c���Z�*@��K\�@C��f����I$W�m1rx��ճ�j8�r����`������[Gj��R�F��P�|����d��$��m�-�P�vEDG�xeM�L�C��9�S���7�M����M��m�)��,���-}X����)�����Y���9R�_�؟ڂ�9���D�=H3˧�}_2f_Q&�оUS�ܣ��CN���K�����57�6��#�M��+�# ��`s�+U.ݵ��'���%��~�Zf�P�c*))��"5Yl�v��A�aޓ9j�L|��}3p߄��mׯ���}< ���4����,y���� �g�ǃ���m�L���<}�9q�7����?��ۺ����+�`&�M�.�~��N݈�S4������:U�2"���������i����Y2�_�l�=������׺0� : �K�m��p��tz�9}�����dNa?h�����f�!'?%���%/��Hk��c��� �Z�j�Awe#�d0g��2{42V���V�èeҰ���`삥�����4���c�֛��q��nEz"I/��K ���]*0ZR�=DN?쾬�t�Q�	77}MX�����W�M��Tzi�x��\��}�i���C['+���G��T0{��NGy90�K�X:��-�{��;�rSczz�ۆ�ȩi�N�d��������dI�d���!H�:i�O?�� ��0u^qq�xO��-?����lk����"CN�сx�$���sհB]I�{b�2h
�]�o�����E  %F"��>f�*~�����\0g���&I���QT!�m�~��ȣ�H�举�X�1@2�=d���L�}^�����1��.��"�i��\�[׻�9��ID؅�F��G��n?b���)뛕G �𩴉�#k�D�[_h��4?�h��XUU�!Ẁ�i�����
p�����K���!���^�9�G��Ui�ΧR�ssD�;J��=+�yM��*�=?~� II�A3�	��H���Q�I���Neݼ#���Y��R��l�	g�G�bF:�98�	�knV:�*�߀H��,��z��쪛]��>Z�Z���H��T-Gmu]Cd�����P�^����u/d�	z#��EEN1����D��"U�Q��
`� ����m�'��K�x\��z��|||ȥbT@Y�ޭ�a}�=�`����'\�8��5M�\#:�O�F$r�距����?-Ƿe�|gݹ�g'!���)��C�4+�*L���%*��n���_C0�頊��2bW�bKϲ~�0^~�V^�3���wU�]����'�˾��^��{��G�f�g.��Up9��L��؝�����q
x�4��89����R���a�~����
�o+���&���]�x�s��	����?�>K�:+Td��G�2?c�hOTN��DtԗL;��'?[-!D����9͉������Q�D0����>i~3$���w_-�EpE�ͮ�J��Z�s�|��A�+��M�k?��r��mȢ z��Q?��fܔ���+]�]Y�:r�'�u����-���4�lx�����H"�n�wK�8�����|�ֿ��ӿ�9��{�w?��b��W4K�ĒsS����ċ 	�!�b9vF��%+�I�����d��M6~������Tྫpk㖇0u��F��Bᠶ�U��ܔ��٥��7t Q�Kư^� ��+�3�m���	,y��� 	Î�N4(���,��ٟ�㓋�4��f���*��tx��4�U����W�@�X�&zBv�o_��/" 5����'�Z�%����jT�zmYXNQȌM���m��V扔%������SJ�JP@�Qnպe�}1�"�jS���K�|�' /4��,+�� �6�sZm�#(�c�(����XL2�
 ��U�[�OW����;�ajP��S�z������Q��@'��5�T7j(ߞ��E�5��qߗ�<C�j**��޳G���)j��g��n`I���8����A�����*��[1��&|g666���6���	|�r��c�V����f��=m�M�t�c�9c�_5!�5IHp�|���
<�ő��y�o�\g
�x��=qf���1;�QCV�X��.�N�iZ����B�Az^�}ȝ,vc�+�>K�+}Qfi�@zUz�pD��󡿓_d-Q���q�\GfU����U�� JxO�;K�)@��;�l.��W'�Vo��g�����/�����	��te�^��Q�l��i��l�Reb��hfjjj��b~�vxҐ��\+����1d�Ć��0}���2�E啎�$]��F�yXfN���v&��gB���h�RZ$sY�}�yal@Ð�Zv�ϝ?�2	]���o^Z�D�B�������-^JWŨ�L#�'������	y "��������Ͻ�E����|<*&�G��H#�{6��V�����J��*犺_�G�g��'��7;������?���?��l%[��t�y�|6lVY�o��b����I���d0sD���=��x\F#�kޢ����a ��>�{��/_�'|"f���W�iP��-�!�(���W�U���nuHj��] &/r97�A9Ч^C��*fb���a����L��-��G���m��-Z�$���M}O0_�ś����;��a���u!h�ץ�"�x�S~�g|��lV�g�%�P��������}����5���h	�b=$����wu����H��L����Ϥ�?e�\\��N��'��6�]��ꄞ�mKPpUt����)w�̴yhmᩞ�"��Od�`Sc%(��D��M�`n��e���9�*�%��������x��z�g�������T�l�8�U�%>,���kd��u��%� ����׾�qF���j>��9�v�Ja�
���m� �qy�ǥ���T̘7��	*"{*�)�rx�W�Q�_e����ݮ�jn����BK2h��z?�w���KR^4i#��+"I����fU��r�NOz�L�)�������o�G)�h��0r�l��/^��J�m���7�+dMÑ�o��_��Y@�I!�^�m����#�6��T��5޼:5��[|��C�df���H��i���$�L�]%]��};����A�`2���g{��o�l�F@�V�Xj~��4�$ee�<Y���_�_D<��	ud^@x�iʲR��D� �IW_�R(��>��EW����Zi��Vk���< �s�H��6��v��({��!-oJ5s��<���x����w�7�F�$%���[��YӊI`,���#����	��~ST�{Sx�#�������S|��W������r"$�L>�������y~�C iY؇�-��q����ɸO`Ζ��W϶[%&Z�b
�e��4��X[ɩ)��J)>̀bI+7.Ay���[���������_��m��CLW:U�������Ɔ�1�+j�o����ܶw�'��b�r&k�'��:�`t�G�uZ�����.(+`�s�C��`���qՖV==�����w�	kȽ�!K���':�$�M���e@0)��;ޱ[����=�)�R�eI�� ����{ �Zl� n�Cb���7`��;�����ӂ	�\��������X�gt�Z��C.��lS�:j�����5��_K�JtDz�9m_�+�mm
Wo�mz��>�W�LJ�b����Y�Y, # ��U�.�/W��6UkM�-U�
t��s��B[�U��8gz��W���nY).�I2��>�A@���sx]%�fm�s�u�noK�r��b(�i�%�����m��<e�9���@����=WE>�Պ��������ϫ\�w(m3�(m��\���܍v�5��&�>j�sJ-L��F�L��_�S�l�C���/r��:	Ft�@���}�(����ً�>�z�D�	 b���2j~k��z��L����ؘG]ޠ�^[�Mc����С��˶Ey���;-M�����;���"=R�����ݔ׹����S04�ß�O*�iTJ�����fMPP��2�'�Qjńk�1<��R�O'J��e��ۃ:��ط���EB�/[%o�%nQ̭����J>O�(��]��}�X�4=-��k���-����4���&b�l�Ό7��z��請sM_З(KV[۲#ˀ)WeJߝ���%�a���S�<�Ѵ����u�$�Y(G��I)�5�5��%�u���뇽��a+e-0R��r���Q�?L��<]v���L��޲�*�p@���	 )�Uf����CV��*2����gD��V�n�৽@���un곮�[�Hu:aIy�T��@�	���S_=[G�v�	�˪���`��'���������$��Ѩ�Fa,ut�������dh!�R[�ņ�|m�5�gV�E�}����NL�c�������H F�1��4��v����ƥ~���8&���,��d�]��O�_���C���nPU=��[���u�p*��3��t���[�"���r���Xt�w[&�I��1	�p���g(�!�b��2���& /@P�X:�'.�����o����ZN����C@jƒ��@��ߜޛ��6��o���d�j|)"����_"���˯����Q#W�c~N�Vi��g�j�rӔ;;9��O���YGvt�o����;����A�I��>���b��PO�|-����؛��T888����Gx�
o2&Fc�:�'^�9�e�ԥ96WZ/V�����^׭��h�[�jxpY��}J���������h.3z���=�������Ό�'���B���l�$o�>�m��ml!L�A��i���M��7F��%�%E���`bП"b:r����aѮ�d���Q�I�.e���5�Ǳ�X�U�N�����{����f���(���-!{��-y�E@�����I'3�b]�;�(]@�gV^^�kd$�椦i�%6�Lݖ�i$�Dp2�|Wj���hW�8[~l��<-H�J[�����F���h�����`��kǞNTS�6����t�� ���o���K��,��K���AT��N �����
�����SǦ�f�g�K i�)HfKb��5�M�D�
Y�Y+$!q%vF^�*���\9�Q�c4���|Z����V���4�E{3�&��գ�HX��	~�*����Z5�75$s�E�6��ϯŁ��q2Qt��7��x)>�[Y��w���w$%����f���6f��	��ÞF6uϒ�� �cE�E���%l�努���J[[Yo}�
�.|gʍl�c�:
�ڳ��]n\c��=C��x���ѽ�{:�w�?
=�U�P�y-V�8DV��hk�-2T���O�x��IF�1B������`��U5����Jv;k�������N���}���[�AG距�(G������x/V�]�DmR&���m,S��fȬ^�#��ރK�����ߥ����5hr��Д�0*6
eRBf� ���L��r����[�u�,�x����O>9X�p�y�-_�kl|���`ð�cǲeZ���%'��Q��=�@�Xߌ|������i��L;�71�0�� �tB���,Y�?��Keב
4�$7�}X�JO#�Z]YzBn����Tooo�`!���U��c���T�ҾCH(����V2�&m�!��}�1�ܫ~�[#(�+���.���	�����?�#wm��`Bt����sL��	#�_zsii��:Q�*��k_K��Z�6�gd�l_]���Q骩���A,K���	��,F�[�S��/�A>~�@�[�ڎckO�3��jJ<eh�`�M�쳱�a�����OK��p |�7�_~O�lXp"�~.]P��
 ����Rr8�DFB����wc�TȽ�j��<@
�	�����U�ȫT-h���D@@72�}�ŧ0Ϳ�n����]օ1ɔב��r��O�����]CC���s-�U�;7o���[	��q�a+��;a4��� �(������/7B#8/Vf���'�H[���?���M���3DO��w�x�i�F
���(�����/>����(0P?B,�ː��h2[�~���>Uƍ�g�-p�BP�����QoU��5����!@�Bpw	����.��]��������o��>�2�cm�{JU���z�\Qb� Ɇ7'����b�����5͊�ߞ�^���I^Vn����R#F �b'~�G���Bi�6Q����'EA��~p ��z�N�ԓ�K��t;�Ƒ0nb0�:>8��������4¡Ohp~����ڀ!����-��nn����QYyoqc����ז�&��C��>}�[C����������!���`:�/��`��o��A�'�/Y9W�R�z;>��`f���cL�Ȭ��TƊ�����������,��:a�?b���=�a�l$�ܷ�3�AP�'��=��f/_��%~/QYGL�QGZ+���,��йO��E�4۲�׾���PP������)��}��y�O�K7n2O���h'Ψ�#�U�vjK��P������� ��O��1N	��H\�V[ۘVK00EE�Ԭ���HYQ��4)���x�9��	,E
�Ͷ&�/�}g-�3�g�X:o0 {#�0`����[��ڻB�ھRdjZ�L�b,�.�{����rY���_t�!�����xs�	���r�Hs�,�����ݕ��ޘ�k��KG?�e�zP���i.�e P��K� R��w�ԁ�"������+2;�wgD��R�ĉ�� t�G�F%6��jZ[G�V`�Z� jS�����mK�� �r�B��΢US^3)0��r#g�	��;���:o�H�^��١�ﵱsX�)�%	n�?�[�,--��� �l|��̙-`�;�N`/@�� XCuƨ�����K�+�g '���\y���V��9WƔA������5I��;xA��eɸ3pI�s�p�C.��w�l0�j~��eQ�6G6�D�oyV��{n���Ȯ�7���)GI�N
j�n2�{H� ���d+��� �F�!s^C��{7Z�B�
b<9�҈f�R�8y�V�0�Mj�:Lӹn١ �P&�3��(c=z���-o��f�)M��ؐƉ3�3�z�(D/��WVN�b�P��p� ����U�Y��Oq����M�Y�lٱ���[��>��������W#��.$��~qE�OǊ�5m+kk&��?�1C1e�׏��g.����CD�c���'ձAo�3�Ȯ6�g�6/��.D�^n�8��u�LB�8'w:'�#���Gw�?e�Ħg��������8�6O�]�s`�ͩJ
8���u�J�6�CG�9��n���%ދ��T���嫦��2����;���WN�+�n
&Θ�:p�f� *E �;�
י��=f�R̦��Xi�O����G��&�s�i�~������:���J4�Ҥ�Js�,�w���ݶogY�o=>>zR4��)�.{Bb�l�"��� ���]��ѣ��=�+YH��2�z��T>���,å)��.9��?0�Bl�pO����%�������:
$Bp_)��_�g��{ hjj����������q}q�eG,��|CMX��ڿ~
�<��Gb�X�zf�_�O-�}75Y;��_dI	b�|�J�On�V�t?zC��\�4kP?/t���{3\�mc��z(y�b�o�����3�7ʋ>Ʈ��2m�]zR��л��Q�}��~ݓ
��Ǟ2O�3gV�ВU�g	���z�;9���@g�S&���yJ�;a��!(+O�7�G�pqY�m+\�]PU͞6��A�<��N�\_�5_�A�

�^��wh�%""��a'f�HR6k�����彵����w��,�x����habL�VxQ��v 'Dc쥛lg�WGk��Kܳu"_X �/"�[v,Om��Jb�J�.�Q������u*��Ѝ���Y���Ig`v�i�5�yo0�FJ�=��"s��TN�>�Q��&5��Qю�X�YȧT�/z驙�%��Ԙ}d��nm��b�T ��22��B?Ű��7��L�ю�l �,r�����
�9��r�;���+R(R�}�;#o_��f�m�z�xh��/q{0����!i�#�l,r�����$�5���P@����*q>��n{J���T�)��>m�w�-[Bf9z�,�q���(U�f��ӟ�#��>WXV:��30%�ڃ��Ρg�
V�3��5��($��OJ{k� (0s�z1	\�,��g����*>.���m�V�o��t���q<R������@����f��Op�TT�Uՙ����nĀ���o����j��O���,��w��n[��O�$ᤔ�TH<���{���9�B��s��=��}�fk�m�Q\�ڭ�G�XW�wܧ�7d��6�=�B�<8��"���}?\��� �K~��pca[Ѿ?�"T��_�۾}M����2U�?J�n��M$���ad�Jh�5�C̐���TFl��,ʘ	��o]gO�wg��Mbޅ�\�{�u�D�Q��o��_x���jRl�G1�=���~��\l�>9c��x.��T����o���ok��6�a�jX�
�A�~�-s��ҧV>H&�W�=T/�!�e�V�1	Ə?�"%`���mT��9-Wm��T͢�����&��]/L�+UN�B���d W�>��Y(�|���?࣓�+�#�y2/��u�3-k����| ݘφ��Ri:^��C�t�Y�Y ���ZL�@����W����}�P�
��t I��uO�������S��Ӂ�u��@g��4%��㻑�¼A 3����/���9��~��E3Y�}gN����J�[8��u�,�%�[��t�䨹����6�d�Y;Wa+���a�h��M�����v4c�㡖k;lĎ}�h�հ��b�ȼ��<��D�.���<Ƈ��އ��Ͼ�2@B݃��,�8MS����'��,���Aw��	XE�w�I��;|..upm_�l���ؤ'62|?C��?`�����uA*�sǤd�gRm��Se���*�{r�'�Yl�,7������6�z]IT$!��h��T^��W|`� t��i_\�o�p�x�q�}Q����؃0e4Xܩ&{0��Դ�f���m-V���=<�6�as�"����BSh�~+����4E�y���<���O���6���[�a�>��o�,^�>�Tv~ܢIS��&�8�v�
����ᦲ[�|I�3����2�i{�4�����V6�/F�8�<f�8�
�_�X��&��+*&r���MI�3��ܜ����DѠ���s>jM����Օ���Y=t%ً��c�cα����Q3�NI�kCq���U�`]H�k( _�r��������۵o�=��AYT�}3Ŋb8y%�Y��ŏ���Ɵ�1WW�1�{o��n��1T��5I-o�{��`�� ��j�D�ՔE�߰���J�;�����S��H�W*=*�6����,"�Om���Z��m0����~L��K�$T�dQv�J��ӑ?��>;J���rD��y��tוr���>�j�����q��;!dDb	���c��ӔW����W�=���Cޮ�|/���t)ת�:E�$�V��v�&��"ZχUKB���'S�˨���$���=�蛷��U~����^D��o^׿��9�b�[����>�_!�_Y��C�~L���`��r(��Ca�a:�ֹ׸�6�~�t �5�Bxjy��>�ಿ�b�8��&�H�M+����Z�[�º����mu��πoWX`��~�|�M�-�	߄����6K����yE����M������m���aU��/��a)s������~�U�|.�;�_�}6���\�G�;��.��?s�~���4[�J����;-6@�D�}{]�|�2�c�\�ⶽc�.c�t#�|��i��d���xk�y�L�#���0��r ���2��a��)WF��cJ<�h�ez'�_v�C���y���%�ە����w�Vϗꎀjߗ�ר5��5��۱�H+�Q��:o|�)Ŝ�^��?R�PJ�HҪ�E��cƂ����u4-5���b��G,�y�7�v����֎H��!-B})�p�w:?��}a�Q�H?�.��R. y���Z�}�������R��\�2sZ�>��Qca��-W��E��@����c�T� r�u+ Г��_�u-�����l �Y ����Q��ϳ�������s���N���s���W��c�&&<��qaW8�\��!��0�G�xQnr��u�_�h]92]��kV�8�k���cR$���>A#�'a{d�!D��IF��4cOZW0�9���o ��-Y%s���ޙ�"�;�He뢔���*��mfy�J�~&���#>�=�!^�{��?�s�v۟@�~Y�k+��`�P��}�6%���}��D[O�	�D�{����5�Ju���0ur�X�/4a�ĩݫ��&-��$L*�ч��J�4me'[nv�=�oB�!�r�.%���_?�C�%��y�x\Q^�ӗ�����Z�:Vq�9�����B��_�������]κ{�K/��߇�uO�'�^_�n]�Lk8l����~b��o���#���<��ı�#F��"���_T��edd&�O]<{���`�J�Gͮ�,����*����G� M��t��%.b �����LF��	�do]���B��$��*�:�͜%�vj&��J��MDq���/��㹿��g����ã�F�Gr�	��5�H©A�(A����9��Kt���^���e�^Nt%�P��''^��A� ��L�T�&���U} �e���Q 2�!f9�e�ш0ZW�Q��\ZZ����h\QY:���|��_ ĩ�ۦ��Q¶�n�,I'*�[��wft�� ��;���f$�rų9��ܜ��0��P����s�Q'��n������0�ʩ+���F�5��\Q���H3 CC�16���5V�CX~v�~!}����0�����׎=yB��e���T�N����z2���a�r�����'�_�ν�T޸�g�ΰCT��'c~����'=h��d�빮i��w����2_�R4��i]�q�����|Uv��C����#7N�7�	�~Fw�
~r�)�?#�q�v��� 	)�T#f�z��#Ưg��t�'ff�"���5�b�YF��*�-,,��eE�����x�qH��D�@�gY��ݼ
�����M_gI����)l6^�8�2�E���R#ij�F��UJ��K+X{�>�~Ι���{�z����n��`uЌu�.[=!��3����IC��1h�b!�n���Ǐ��!0�#�Eеv��tc�~�[Ï���G{B��l�k�'L~��"�����S���!�³.w/!�<����k<�ˣl�2P��~����r�� ����I&�麍]#c�n�HQ�	k+6�u{Q1��蹳��a$p���Ttd��NN��,��$�?��fg1�+�b��ЁA~�l�\�� �:�����-�(Z�Q���v#&���̩a�[P���o*�KAY��.V"L�$4$k��/:�¯�2�i*�\6e�Ѯ��7�`�K��άÓ���!{5�n�l�蓅��֨�ţ+�_Ӥ�xGyF���苊���A��q�ef���a5�3�ͧ� �`er�	?�ϲ�)ϰ�8(�B�1K���L�F�Z�5N�k�(ёNG�A*�����G��S�M	D��<g�oN���	ůq(E-��C�:m棰Ӝ>��
���[�N�,��8��� 3����-���ܶ�u���l`�&����q=��~ѕ�2l\�+N�ps߿�0r����^8�l�>`O8frm�I��s�=}�
%����7�B��sگ�KFˢ�Y��Ҕ��s���A:�|>هNm;|h�o���r�&�K;���eRRR�bKHv� �WCs�����l2�t�рw� ?໔h��I��X�J-�lm��%5+nno���`���&?t�&�گ^y~�w�?-����q��5��Z���d�+�WI�&�p�' vy]�����X1����YaCq��:�>���ȥ7v{=m�gп�J���)h3�j�A��/����9A7xQ�n<z�j�#�H��v�78���K�)[�\��1�&�G������Þ�<F4I�#�I���X�v�z��0�� �:����K�Ș�ry���ň��	����(m����-���o����Rd}'�D�=���W�5�[\+�B�u�Uޜ9�	Tt�NMd�Dcc� ��w����NS�@�'w�!n��^�����J�D@_���p�L2�IC{o v&���w�M����������G�J
K��5��!:�8y�m�YP*-�2�}o�s�y�E��bv�Ņ�	5���X'��R�uK�ʹ�^K����$WyW�t���B��n���q�AH�Z��e�0��$IA�X�&�}���<���K}��8��8E$��6@e6FΡ�dq����C�C���|F����`8��J:�t�e�/���τcГ����D�D啵��h��d��{���@8�b����|�H�m2	33D�Zt�-9�13���K|r܇����gw�H �*)/�����$̋���#������ztP�V uppP|4+zGN^���o���'���kn-z�Xpph���9:Ď=rkKvv�E۪��]�s���$=�E�^b�!a
� .FFF�~�/�^YA,�++��0b����3��}�&��MWd���"�3VV֞�{C3��]D���%#������0 `rH7�=mָ��k��l?.H$����(,h��(��}�g�*Q�M�9-�S?b�;m��-Y�cj�$g�P�!����ðy��!�Ղ$
�K*��p;��e7 �TZ�'�C�T�O�?=�V�o�"�Z�Ch�Nw���Ay��{Î4����d�3Z�v�b"2����i�WՆn��Q�9=�b�t�-��L~�-?������G� �����w�H�E�B^$X�"5T��N&��Dɑ5�ћRUE��؈��^����Sv�ԨFkfe4gA��
0L �D�	U�.��D�VV"E��Ơ�9����pa���J*+�'q����	������LM�#!!�0�x�遱e�L&b F�y'�7<�''[.R��x>R&�����JTW7��ex���e��������\�7�8���̨�!D\>M^�TWW�+���s\��ϕ˫RM�j�'y���Zp��i�����̲�}�����tu���e�͡����xO�.���b���-E���m�GH���]�`��h���T3�m]+��J����1e�BS�n-�3sn����Z���1Ғ>�j[��ˎ��|����3���D�W�7DZ�����4�N�`�7����4ҫm�_�<��\�e��p���x�j���EnW+^��4��rL�������(Cw�A�'�ۖn���)���G��52M�`�2�7�*���%%%rܣ�ff�]��ش���_�K�BQ�E����v� ���h���ЪCD���dG,������qA�PR���^Iu�*���=hjf��^ =�"~���=:���� �$������Y`�	 ��W�U������R��`/�y�@c�
�N��maάA.�N����m���
�Y�E��Rjo/�_�����ή<�*�o���`~�����Zq֑�H�v��G�T�N�]$��oe�����ػ�q���j>�9��nIS�u������09��!SAI4����k̤�k��Uj$��kOǙ���_7b/��/U�dy���Dc.����;#5G���Ci�
�z���J��?�I�3�Yː�Nn=hu����(�Q�fg�����vw���I)�{ܔ���4X[[S���?�^'�4nŒ�M�!8+�U��l\k�%���ky�ʞC^eee	� ).R~AA�ZQ��NO��k�j���î��9�����хg%���\�OF�r�[�Q�B I�$!��6ӣc���jS��^������49i�TiPq!�_~�c����9�a$�IS�C��l~H[�X|�� �u�0'����ŲC�WB{�k�㠇���ν�rވ��>����x�&\��aEkv�W��&>쫰w=�]�^ь��6$��3�d}���U姜^��̏9��Z�{I��H� w���;b�r����]}mm�P)y�G�4%���KmlȀ�PL��O���%��r#�E%R26��V����?��	�^)���1�����'Rj1QQ%<�w"�d����r�:1ER)}GN�N낗���;��)�_�$��v�ѕ����%��\[��ڜ̧�W�` ��J466�d:� :�O�>)���7�!�1�::L��_��dq�e7�g�iN����b�l�m��{�����R�Ŷ��G����A!N��� �z��ͭ�������H��T-�~��ύ����ƌ0�R�SP+29bU�zoo�$�;NvX�v^�\��/����y��_]Jv��p�.���v�)�	��+�Z��<:�rM,C��|�{p3��E�O��Vct=�0"�:������eW�|q �z�a���m��/�r ��������CCx@�y8Upx��D¡
����/,��qr��ފ���Wa_����2�j��b�/_ߖ��~�0)�~4g��.\ɴ�c+���_'���)�1v��x�x��=_?��'
b��ǎ�'�W����Q�v��H�+�j7��1m��[�zQÄ\�C�8�%�dI[�7�a/����]�82�IGX�%�BO^��,����jG_��%~���6Rw]���p��r�޿<"�)��惖F'Og���:�̸L���R�-vӸɗ�>ʄ���vM�+y���!aQJ�9,��+~�(L9�����x "s� ���?A�z!��i��0!|�L%8z���;�t�	
�t94,�x!﷓��z������=̉ ��P(J^y�T�սg*��Na%��Vj��MM��,i�f��q֮�c܎�����.�h �u���\��R�i����V=	��EV%�,��*�!�N�J=m���4�;���,�0ͫ��~��|���/�q��	ackX��4nċУ�|yj�޵[8}����:W��X�/`�ݐZK?U��ok��"��^	j�).���hʤ ��K�s*�x��]�6�c�ȴ>[F���~�J�fl�t�cqq�Y�  ���AwgB��bN���c���S�
�hB�:�;/�9<;x}m]?�c��R&��������$���d%jX�3����ٖV �@�����h�e����	�ڝ.2)������?�yIA�֩5����\���!�y>���7q�&#$$���� �j%���Ed:��05P�@b��b�8�|2?���Q����GL�3�0:��Y���D3�����P�	ڃ2�hA�0��=Eҗ�h�ϧ���A��5��BrL��"UһKۑ�j=�͗�O���-A�z/�=�X�����C)]�ڣ
Po�n?�+�g:)���7��)z�~w�V�(P6����k�{����]�[X�ה����u*�ȟ���i�d_"\�ʔ�/ohkk3Yt�+i�i��HdT��� �.ݸ
舀P3V���Б�)m��:��(� �d����m�ch����O�:t�$xhg�dœ&�D���DpPeH����Mf�� Fnٵl^��^�^��h���ժ��T-N�1TMaa��I������r�q& ����o��K,P;!��[�����+������u��9����k�QQQe'�::�z�ԥ�+�(76NÿT�v�h+kS<��0���Q������V�%�2�.��s�+O��u��g�Yg�I^�{��Ѣy�7pW�I���a��$/��@���(b��q�@�����|���9b�Z���7Tj��L�5��;HƟϯ!���bz\���]ˮb���4(7��мe}/+�=�=G�>#漶�������H��+M[C|�������F��>$h�$h``j�*� `\$;B���pR �+�bn_����a$c[b��m��V5|yY��s0��ic7yy������M�{j{�X� �hG
$%i��W��P�<���cvv���f�-P���qd�E����]P\kR����ˌ5��1����	����C�pe�iq_]�)�~�R��/A�N����88` ��~Wh)q��_G%�ߝE�o-'� �P����c�#T�9�!!0P��ݕ*��4�MMl�:j�ܗ�1з��g_� �<@z���[�uN��W~�=�a�M:V�]���m��*����.���I]n=�&�B�s���{��y]p�A���n�&R��^�t�i��S�ۿ`'^qB�t�R�^ߝl=lO2^vn�����B)5���uN��?AVC��n��`��5�@��M��4%���x`�FiI���-�	�	��u��م���6���v:�0 �a
3�qg�s�0�G�i'��`��I�ĩ�R�5��VU���K'�4�o�ޫ�ֻ�,�ˍ�H���G����ς�[~�����t�;���ͣ��Ч�d��А���=X{����Kak�m��;~7*yp�ǉ\�aK��	wL���J�8w�����Z*b���?L*�Z|��ݱ�&:� 	u��O�i��	߮*�?XM�q��l{!��o?y{ɞ8�6u��9z'|���l����t�Uf^#��
��L�s�M�ֿO�
�Eee������>��/͗/��?t���W�k��On�^y��噊s]>����ln��_�*�������=��vjۉЯWM����-�*?@��8�+���o�w9v-[����0���(�b��A���S��bL�z�B�m W�e�c�5�B�ǎ)Ņm�)�b��2�ꋂ>Ϟݚ�7���W���O>1A�u#@�qO�N�<����c�j;+��z��Uq�ZėpX>
7�;��]wX$d�ȿlOy����j����~�k����J;���Z[�i�oz�B�2gCf<"������F)t��I_�S���u���O3����2�=܂+U�	�z�0UL��}�,�,=���]ç۔8<��XZă_v����}��@����ވ��߮�5<��C){���V;$מ�k����8b��t�8 ��;.�2W��|E�g�*���J�,P7���Mc�]�P�Ȩ;���~T��ȝ �b�mz��_�N���`�@8k�y��w8��Rc��z��n'�Ɓ�W@۰�wA�z�T�#ʇ`��e��yd!m	����e�nAڔlv�i;���ڔx� V�è��!9x�/3��j=؄���}a&F����j
��I��f�-����5Ʃ`*�ڹ��B�����19�wϡt��q�.]�0�֍�h�gE�4K�5|�RE?��i�ّ�#�L�uf�Ƹ&�Rth<�6��mi�I�8�r��^nq���)~Uo�,��3�-)�����;V�K��0`;[}@�w��0��	��r|����,x�����f��]d_�Kf3ĝ�
���W����
[�ˆ�j��0���Z��o�Fp>��E�₼���{�L�������k����?ߋ�#'S�5~�~�E���r'�F\j���d��$�l|�����%{wڲy�Z���o���su�å`��DX��<{��5�'�?'�w2������@��E�&/Y��~R��Kv.߰�FR���C3F}��.+,�̯Vm�yU*��[��A��
���\Y�y0� ���۳/��/)]��<��Q@�5ō��<�Z��"S�����]�5{��;2��5w$n�9L�=�|����~~EĐ�yMU��OuDE������6|����/�c���߯�����5����?����Hc	c���C\c/x�+&����e2]rW�����]/�1�h�x�4�nЃ���Z�p��H�|�~�yٓIm��=-o&6(��hR�ת�g��nfu�~���*YO�����:S����' +�%�!��ݑ@���������W�ar'jr̫��R�
�<ߛ{w
j��^F������&/��P=Z��W��.�-1ĴЋ81W�7��,Z�4-=5��UF�����Q�M��dO}F�}�q!ce
Q1Qc���x�?���qqq��S'�5j�a��B�zt�|@F�%/���}a!+z0��1S���R ֭~I�B8bct��D�)W��R��w��;�̸�/��镙'V��	�k�
�0�߅λ�$��08<b,��~��E�14�8&�~�(�"����j����T/�!;��^��u�E���v��p���DW{��M��ۮ��F5@!��J���_�M�zv��������LT[�ٿ�������U��JVi�:M�3�y11L��:�>9�l�NK@��[�>��@�ѴIU��<����l��Zr��@	���t�_�'�V�V��s�`3�D�O�r���	V���|M�լ:>ƫ'k3�S��i�
�x�R�h��*�l�G��u�҆.rQC�_�u�YU~�B��>���9��X�VÃ��w�=�	A��
j9k�A�>�C��m��qc���8���.R��@.1$Bd�����7���7݉q�+HFHъ���MLJ2�`����n��0c�)6np���X�px�!��w䮠���!��.��`�x��|*��+� )7וǜZ[B~&�d�����
,^bK����a�����W�����j�ӖxD?����:Q�!�g��=X�ӈ�ar��Qe��מ���^�HJ5�WU����۝o	��y�r�/J-�4�m�]�"Y�S��r(�t��}��[
�]�J+GZw���;���MOw�uu�������ڠس������,{��Z��!�ac�Yc<�g��jl�X����lm�He�+{�8uPx�/��6�yX6]a}rkd,)�T!t�`�y��d>{���Ȝ�e;�|�U훼�+��An�+S���L\���_���L/��c����z?��1�Ǎ\��7�=��yD8T�B�<�I���x���������Lh��"�+��i\5���� 6/ ^(,�b|~+���iT���u:���d×�a0X��)وA��v���K���þJ��39\�|�l
��_M娋0�_��-��^�|ޫ��?��Y{cis����o�Tw�Vl�H�R��"���3�T��;� g�:��f��y����{"5�_�T�u� �t=�mV�iS����oG��q�^�s�ht,����oO=�8��$�;-	W�`�G&�J�{)���ީQݸB�DW�r��w�Q�!�0>���ɶ4���,l��<a�v�Ԋ�Ox�G�l 
��R__l5��\a{�kV/�E��f�^��]q0��y@Mh�p��g�ϭT�OS�zZ�LV�^�~��=�Q��޾����O�J�u�?�
�{��F�`?O��l�U��3x9�e��Ϣq�)�`��/�crQQE�f�UoAo�# �h(8��J���	LuG��پ���?hƞ���cӥg����b�ԑ�<uѲb#(�,��qvv���%qA'�
�:�U����"hi��T}�.o�J����2�&3}%���pcZIs���zG:g��z.*�Ϟ�����K����m�*Y�w��dw��	����x0�a���X��-�j��~�C����C��.RS��՜���o����uG�4�M���mєmu]ʟgr��[��o��!�҆4�������+��@TU,e�J1e:f�Ls�x���j��}+
1�?�H�CpʢF�\��2`�Rd\C�|H���1<9�y�`���ѳƅ>�ă�����'$f�~|`�;ݐ�����]�/!B�����5E��X��{�}��G����J8������a�>��j�eb9�l�)�y��ϓ��x]��s�Ћ��a$dL��S\z5T0F[PM�5[��vJ9zDQ��d��ޛ�D\=�m���vSJ�%��}?r��A�VX4���Oq�lC�p{�+7��ꄿ���%G�O?d����b����5��5��z��#?s9� �i�^�F��0��<s��d����SAA�cm�f3
22r݁�\7�I��tW�4�#1؊�zbe0k�*4#�h!�G��O�����[	���\��l�G��x�j�����l�=],)JȠ�V��ݻ<�8��F� �L���MIh~Zjü���w?q����
�>?���¿�P��ڒ>���؎��=��C�SZ}�&�"^��p�Rǎ��{{�{�8�d�}9ꁾYw�;�~]ۜ]����ؿ�X�P}٫j�M��y���c,'E�0Ed`�"�q������KFN�yd%#�'���#��3���jk�-��xr B$c��������`��1v5�ֆ�J{�}�ke����Ɗc�QBU��ke�����0k�l��n��<K�'կ���T6��Ä��o�q�>�Ë�� ��k�A0F$B�Ǫ|D��Z}�׽hd��0���_ޘ]-�9�r�]��x?9ּ�t�������~x�Z��El��@f���~�b�[���ns�\���}S��Սq>��[������6'U<���3�c<�m@g�(������� ���X��ӸV�b)fHh�5}G�4���Yc���Z���6��Tq �G�`P�X�}��t>vlF+f����VQ����`x�?hfo�Ic3a�n�bl8%������R�Âb3��j�/rU�Ѭ*�<����p��D�sD����"����h���xڣ
�!ԉ�}ɭ��W9�Ԝ!���\����[Ԡ ��[J2(Z����a�Y�#�����o�:c�G�*P`c_���n+��لgZ6U���7~�ESL�
�����|���j��z�~F�Y,ACE2iʄBoh~S1�H�,����Vt�n=YN�˅ݱ%`Q��G_�'&��=ZL�U>�oB�;h�o6H��3�i������_���Z�a��r;�u�4|"�J��=a����u��H��Y2��W;,��n��򒐓��^N��"9�k�QW�5�G�'���5w@S�,G��G��N����(**R��wo�j��R��k�JP&� �lov������N�?4$�̆�����`�c4���*���V�c����1�$
!@���N6�����E�,(h@��$�y��[�����ŊQ��փQ��D܄��a6)�ܒo�79�B���Q��Wڲ4D��~��r饂�:�:�WQ8���r�@���1��G=�1��Ȑ���	����0�;���9�Y��j�U�����st�*���P�#{��b�@�;8�7�ef�A�V&H�b�����ɹ|�}�@���'��Ԥ���3-Ő�C<y�6K���f!�jM����Z3&��Ȯ9h����LH0y�����DY@`�� tS�����#3, �Ocva6�	`콗�mo�*��cm�O��b1)d��5��.S��u�6�ĸ���bxT�ޘ��_jL0?�,����L��D�c��� �SVtoz=c�-`Y0��봯D'0�A� �����=@����r2���~�����y����f'�v?:�?�U��Qr�����$M:>9G�����9�1L%ڛ3Y>N�H)c���'���C����(Q-ߗ[wJ��OH0����'�S�7��}1�n/�l�D΋�?��}.���vLC���u
��e��櫃�	N����W�?��Ň�`$W��h?Mlh�(F{���?=PŹ���fG=��=l�Pd)��R�y��vA|"�������Z��s�W��)�/�w�O�ktÿ�

<�J^/��x���t}��4�Z<��n�q~~/����J��h>�����9AX;��G��b�?����i-���=�FP�lV[�!!!��:1����{p=ޞ{qy�HCC���&�<aD�.Tl`Q����<���A�$I$>��WnZu8Υ����i����>��XI]]��M���Nܧ�=�����-|�y/W�YŤ�'4_�Z����:��`�oZ�JA�%�ƅ���z�q�:1�vğ�(DM�MF�Nҭ��e�����85T@�8��.8���?�:>U%�ŧ}Aa��?7�Dj�d�L�����v(!�x_�8L2�?�F�����G��S&�����Mm�����{=E����P�=�3�<������Д�Cwu���>�����a��?sK�H�s�!�0Kj��ڰ�<��ߋ3Rd� �L���Ee5�f��#&VuNn��%��MF�0���k��$sK�#L�>���@O/7w��z��x4�.�'g��W�ȴ�Ж�P��{A&�֚�
��2�*��|<������nQ�6(�	������	�G߿��C��l������> l߹�ԃY�%�7O�j��{d�J��jLP��m3�H;"�g9�'�\�g��ځ�oD1�(&��Vh}�!���=�b�"b@����
B��\<��&a.�O��H���r������b9����E���# ��BP��T�+*qz���'�ˋ.1���Hk������U~���s��7�V��Es��Ǐe����Ek���~ɍ*�F?B���_�	�o���yv˥�B��Z�9���0�9t/# 0N]��LX"Eɜ8?�GC���w�89�	&M�m~=<;��B4�\l��U�M�c�57�p��i���
�1�1��^�+շ�طe7a��q	zIMOW��.����62b�f:`�?eԫ��C���4̈ƕ�����@��Ӧ����W&&p�����C!���DT}�H���M�#F�f|�(kz�Z���4c4>��q2=a�|���`4��f���e�V�0�Y\;َ;Ҡ�"s�VF/=d�f��j;���j�X���Xٿ_�	ұ�`��v�MgWӴ��	n��]C����.�	�\�;w����-Ȣ�������y���ujY�=�w_=�3���W
����v�@���c��.��ɜ�;%{�/F��ۺ�O�%�OR�� m)�5;��B��k_�ZwH:�|���g�3�'�?��c˂�'�����ݾ�s����"��e�(��nSlЪq�JZcq���*%�csY�;BN۞j���%��������9X����'�6�����P0�mq7D��� %%�Ϻ�2r<�Tp�#�G!;�h�$�+��y�CN��h^�$n��;;l�bu�(�#����'(n�[	.o
����|��e����]��7���g	H)v� ~++����7����C������������G����M���l`�7�8�F���	�R�h;$�D�����30\�w|�����)au)n"I��Ѳ}�g�Uׅ��-��u��L }G�[�2HJ6�!���FO 5&;�Ⱦ����i ]�)s՟�F�8�n7SƦv�Q�&�τ��s+tX؎��$����u}�T}5b�wʗ����$�+Q���\�t���[��n�!4��-(S�G	5H�vogdLv�A�{�ώ��e�����Z:ʫ�T N�F��ߑP��}@�B��"*����*aL/ [��$W\M[�)�M�֜@~�k��y����s��?:ꏧ�r�O��BB�w&
��pNJM���Rڵ�J: (������Q���P�N��6e55����E��E[ITv���o-�����J,-/k���;���d��T���%|�6�������h��aG���k�b��kt�}aMW��EN�P�I�,��?77�&"R���ߧ������*:6v��ì[5�" eT�B���������`��m�C}�a@6�������R2�����T�A����U���ڡ�p����L����FO��eVxJ�#���C����2Ii
��U$�9�K��I�������Y���y	�u��lՃ��|�_�ʧ�S���KϠcP��-��n��u�du�e��Q"` �<��~t�n�9drhVK(�ϗ�i#���a�C�W������U.�$6L&�A_w2n���^������������Z�o�5��3���#'gŤ����R$@p4ڞ��@�%�����Zg�ΨS������cھzF`xjM�Ե� H�4��ӅR �I��@��W��BB��4���<.j�镕�Hj�u�݊	 ([{$Q�S������b�������c7�c�I=&������)�1[���Ĺ�֒�򺻻���3�
��Tn��AeE��6ae%�Z9�URǥ�'$��)߄ۼW�H����b�1��{��c'����~����(}�Jٶ�Q���G]�Zר�M���'B���2P�J3�����x�ΰ�u�z�Nb��32�������q�*�����]��ܿ-�Bq%�B~�4�^�ܨ���8/����裲L�U��!���]���c1v�ο��b�*�S(�0��/"N�[,���{�%3��saA4��������
�^{M��Ç���!"2,h\� [��o��Up��:�111�VV*�́�&��fe-������|��g<���$�? �Qpvvv���?����Vj׉&G������B=އ'�	()�/�V�^��<��Z���BP��������W�ͧ�l��U6�tʐ]y�>�GL z6�� W]��a2G�q�=�g�r�CA�1��)��V㌗@I.�y�����=���e
�y���
~+:TQ:,�f�������o,s�׮��b��Y#n+�.��CE������Z;:���/��X�f�}�7�g��� �*�p:"��6�� k�>��������l(A�~I�sq�2����k�֓�"đ;:��k�	EAg��B}�ګ��)���j�`xK;;	�Q���#ʔ��!��3c�%6O���҃k/F�f�����ޘ�0�T�_K�ҼG{���vV��8�8��pn}�J�Jޫ�+�G�뢏���р :�����?�� *�q�" d�t�rws.Zf����;��ӆ�`}�B��v[��N2Kֳ{�)��d_/xu�g�F�KVܪ�\�Y���6�MP�S~4v+�B	Qu����p�3����0� p���g	�r���?;����zE�&	����[�O�����jK��K���,(AQ�Ɍ�^��_F�i94�����XF��'��W�V��&�$�9lĔ�~E����]�PՈ�G�02"nG��ޛ�r��P�)@W2�l�w �s��ԝ�7nr����em��a1�о5��=Zjj­��������g�E��@�h��bh��������;����_�/TVĠur����N����@z��,�F�b� nf���%$��C�f0�X�4y�ˡӘ��Dy
�u̷ʔu����|o���D�ua/6��e�
�ňJ�v\ �<[�%T��ގy,+���%KIp�[/֨�L������5������`��%� �iq���'- �:���\+ҽ�)
�YsV��T����m�a��ӡ����-�%3����%��'������kq�ٹ��r7\���娛7	\���	RxM�>��|:ί�.*x��(]*�������o�X��_>7�|̏�Ɨ���הu�'OږRVQ�g�R~�Yѿ�o��	<�r�Lhf�Q��>���j!�d�wr/z�r�D����� a]ك��+�� �ݛ�&�S�%��#	k�D�%�9
iϯ˧�	5v����KZ$��D��ߺ�R���}P�$�o�He�"�Ū��CT_�2ni_h�1������10v��_���-	��#�uA���/��4���Ka�5"�s|<�������/_TW8-"���T�����gT(6DTT�"3PZ[uY�5|�N�b�)�A�͖	�4�����/7�t[p�eX����~N-,�M�┟<�o-}���ro��>���3�?%�
�a�3�G�9d��>:�w^	 }����n"U1����s�k�bl�;ԋ���3mO���Fo<��R��R ��/�ň\�e�g�IC���P~�O�K����EMt�?�a&}�3d4��`t��m���s6������Ї��8��M��ɛus���U��}�.�_EfDa[��ٸ�0�]isK�VO ��0�=�M �C'ej�׳���2�d#dJ�K�ӡ��ƣk5c��!`������E+��g�W\��X���+;��:�-6  �^�k	+"���/�}ĳ�t9��t�G�{��"]��EMML@xt_bd-����Y�ÝG�E�[�3<Ȩ��g�2w���5������z2�}�b��'v�Ϣ�c�y)�6�}�k!%��:�������%���֥W�f,H���9��2^b�w<�w��H!�~�q'�F�fj�rmJ;�����6s=ND@�R�5@ap,��U$�����h���[J0�.�s�*���B~w7�����	0�,$�Pԍ��"�����%�pF�d���~�5vq���d?��/m��C����v����Zu+\��S*�� �x�d �����ތ
<(�<?d��� b 8q���߿5�57�V�֪�݂���U��	��I
���zo����Ĕ������-Ϣ��k+�?�5����I��W�4����)SG:�Z6�?
��ݒ�.☽���8i�������7iͿ�H�_�]2����T�AS{<-�Xq����Xh"�h�=H�2�U���6���:�z�De��R4	�F�%׌��
?���d��V1�Qfb*�6X�������l����5������FX�Q�� ��g�+�#�e��e�-^���qk9��sZa�mē���� �!�|O[�p����%x�EN��@�dd������aA��F�����i7o�txx��GQ�׏�ۀɧߪ����=NԡƱ���_2GL��4���!#�v+�?���fs�3]�����b��d4[�B�~�BP�.{p=��־�";颉��;v�j�f�+B<���vK��������v��QRwZ�p�|���[���5�m�/�-�}GS4��S�3���?)�p� �?B�k��Ur^gt�ڗN؁D˽�zK/�?�5^x�P|!\���Ҕ}��чjD<z��]�c�K^��L�E�$uKskT��E�:�C�.#x�H�n^i���()wb'��'7L4����;̾�x��{�y���rj;7*�V��(��t�nDC2�:::eK��zE3Vo'n��y!���W�_����@ޚC�V���"��$Ⴠ+\�"|h+�F�D˻+83����i3�JS9?�GHf���O^��ʚ���q=钙�m�a�C���A���������朙�uq��t�ʌ��߃_l��7��|�����\�\��%
k@��qGֿ��:��i�����?��>���2�W��������,�J�yí�k��%Z_������ԇ��]�赡�p�&���-�G3�w��&˷ч����g��er�J�\&�{\�4~��[���h�&��8����^\�L� S�|ݞK��%j!URY��w���?U��Db�X;E���5k�,�ѵaA@p9�p���n蘻v�F���G��1��kBb���3�"3���[o-�7���h����~����dOW��¦gVa���R��
d*Ji���5p-��k���?)��M��l��W�����TW����^'���*��~�g����1��A�h� <�.�i���{�g"�&�l��T�\Է��s��r��q��<�����i��Z��}^����8���g���W�E?��^�����m�3�a��m��o�ߓc+y�m�\�m�X9CD�I�ɓ���i~Ѳ��Sx�nպܫ��X� ����2��gS0< �_s���K�?����y���20�oXzIn�{���P ��QD��xA\UYI�1��������EoO ���V�U��y	������E �9��c�Oڼ�5�Z��9��z�$t�7��'�����%��<Z�s��H�T^� I�x`���H��Z�"L�}-d�[�w�g���2�~:����p��{O���˲�B/��~��]>�C!�e�����#��tI�w���ty
�  ��8~��?tM���j�%^�՘���e1h�z۲��0`�����)��zΐ�mw�k_��$H��`����<+����W���		����F�5Օ�ؾu>)y���[f%��������G��l@�O#��5�֗���7�t�#�j3^�0��������~��R����+/$����;��c�U�Z�Ͻ#ե%�����j���9���#����ӗ��ӄyUF�n+���ɤ���#I�e�[�&�"V�#����:�Xn�:�ٌC'벑Z��en�}}K�n�Yru�A�&'�o�Z��QO�U��P �m#��"���yޯ���C�G)��Ǔ}.��~�o���9�u�5��gl��h:K��G����̯�j+Cd�jh̧Z�"���o]5E�>%	�p]ur�m�U˒�����ԣ���c���Z|���TX����Ǭ�D�6դ��z���C�p��k҅�z	�7mUst�����,��_�i�Ts��E֥	M	�^������zn�i�HY�����s§X]~Bz��r�i��V��&S�
fX�\�7�nA�rק��[)b�:&9,�wS�eo���n��P�����{k���p�=������~���?<a��k��^��>�=�j�6�n�h��e۷K��-�?Ny،�7�A�8�����z"�<�.\W��t4�s�I�*z�ë=SuOn9|g�vё��g��Vy+��u�w3e���G<�1D��A�/�i�ڎ�B�)	.����S9דD�}%���f���[����yI��M��?$K�2<x�9�b����<��Q�&8U��*�\����	=1o�p-}^f���V��4��9jS�f>���O���s ߹�2m9��=	��,'�}�Œ.�s��ΐ\_C)H�.OS&&-W�WN�FM6F����iZ3=q�{�c�L�zb�&���4����s�m� �0놽�W<?�+8���\��e�����r�������S|}�3I�J�߾�G�y������"3��]�*�b]��Td�bnoñ`�Փ��z�.{RS&ڢU�v��Zk:��%9[��%:����� �\�0�wz�	=_�6!ǖ��]������~6s5��!�7�Ⱦn��iT�I*M-�;r�Ӷ�9hE���9��K�XrJ��臚��F�~�3�N ���@.}dG`"�:r�Rv�0$s=���65���m��Wb��'�31���җ�'h����,M8��Y��g�/��i�m���i�!���c�y~�]���~��^5,1V������;kc!�K����cE5,�n8��� ����)�84ǟag�F\��Cyy�e�Uh�+O&��Ȭ�!DԳ1��k�c���
��������,_���2�H3��<=W����$gV�$ӝ��h�T�3��kO�^��n���.�ɲT�?�-4�����|��~��6|�3t�I���v��g2�&_����I���D�=p����͈[i�-X��VF��9h\��1�,���Xf��!|p'���/鎽����`���̏���ŗ'�ySmu���O��:-����N�g��K���������nQ�Y(�bk�s��Yy�#��?�m�>��.�wڅ:Y����?��3?�D�}���I����Ez�f�3�'�<�{��x;����Y�؉Qa�_r�c5]7$P��W�mi�����.BTwL.(Sw6��/�=�_��?yfG-�1A��6筛�����ZO~�oNB&�
�Fn\n{����'o�n[�8r�97�@QfT�*u����$[V_ީ}�z����>��p���.C��W�X]b��z2���2�lޟ�@��]�C�c��<q>��Fޙz��wC��%�;��W<x⟴@S�A��j2��MȗL��s�����/)��%���t֚�����85������y�~�X"0����Y��M�b�K��&&����8wb���o{�ڳ^i���d��S�����^�n�tQ��V��v�� ��<6.�N�4x���� ����T3f�MW�kߪ <���VGwI�]6^��Ƈe.=:W~P������{C��$_�r͑��� ��t��������{F,1ά ��� K���\�$'�>�heF�[J�����cd:���ӷkXv��/3���_5ϷY�5�;VBa5zЏ_&������̽K�s�UÄU�IN/���1ۧ�s%)3WC�/X)�>�E1w�!)�~߷��cc)b&������s�_5�����_� ����;�*s,���̻�$G�UbVV�����\3�N~ݤ���S��p���7�yI��}{�	[֟�������n}��L��b�/�@�S��x����j�e��L��C�Y���gJ�8s8E�'o}M�G��6DPesCҰV��'Ó��ZDI	:LÖ �XC���c��M�6V{U-
x/�R�H KD,k70r=�#C��7��{K^]q$���\� ��&>�bAb�1?Kq�B��7M��o�+�xSZ��}bgw���-���RHY ��>X�Zf�9iPϑ=���H�3��'�'3Fr��
�_޽?h�h��4׌�G���(�A�|}uQ%����
�昳�wP8�W�V�4;���^_RIkЯ瘻�-��
&�i]�r��҉�za�����ِ�=���3d\������Ht�_TN�ҏ����"��=�7�3����eد�ތV�����L��ɇ����R�I@�<�V��^�,��������g9cx: P�ڧ�D��߽�t?xy{�Y ��5�Y҇��mx�h黾5��3Y���7h"����(MU�f���q��U��i:V��!	�7�eHF2��>>��~iEM�bI�%�ܪb�O8���ں�X�fqS�>��Db̗�Q�����w:L��9�ޕL�5�[�l��7l���F�Z��N���^+��$�a�Y�1l�����*�����5,b�V#��ȡr,#���`��A�up���`�m��O{��Wsj|�Y�k3i�ݟ��v�bhf&�:G(A�7_�.S#�x^v9k��Y��.��E�Q�#�ဒ,	s�qR�Č�n�q������~N�UQ�q?~��l̃�"
���:ٖO�/�)��x�@4�:+S7y~����caee=Z���cb
��>(��8Y��۹�C��`R�=���� �sx�q�5Y�L�����uB�,W��/���k����Ǣӹ'a&�Yʦ�Z�+���(���eEhf����qzT%1�!qr��ʖ��#]���J�7K�Sy2
���wj�'֯d�M��ތ���<IKS�!Ԩ��I�jNS��Ŀ��7� \*��O���1�IUB�{��/u*.9�x0r�������(�=$��;:b�a�z��b��%S0Q��S�jFy�ۙU�!�B���P��1잶������|�nY�!�<E@��io���3{�e�W��9{*�a����u�^���5�q�>�{c�M? ���e��D�ڇ�q�M��2��6β�n��2efy���}�껨���+�	n��/��6�(��w���Oѱ�}�}�S�'�8�O)���At'$=	i��rĲ������@�AO�A�$�7���{h��;K�s�1N`�u,?��fz�x�������w��R>�=4�	�����E���-7�+���F�7�ȯaӇF/�i���Y闈~8�j'ՕHX��3( �9C�n���K�-*rwڭ{�BɋĴ/���P�^���ԡT�
o%�tΚ�Ѧp�p*�IJN���7�1���"�pѢ�9{|ƟT*V�����R�ɈA�,־k���q�E���ER�jY���s��b��E����S�O�h�F�Ж���B ���K"����v�z'�.;�ڳ�\̄�$2g!�ag�u��k�l�� ���ˠd{����s����ڌ�y�_�������b���l�lZץ�V
�̭��jӛ���԰O����o�+㿥՛�!K,9��toLE�-����K�l �QA1�����΅����HuI!)q$8������ώ衭�Eޞ60�S��WD��ɽD��Ɲ7�,�e
�*����4����>����\�!c�)Կ����Etq.���]}y	։W)��w!r���M��3MY�pƔ�$���7��y�0k�P|�^�g�t�C��0�Ňv"e��o��b��3Ί-0��&�;��ad������a��	/�j^aQ�I�/��C^��ƵFF��^��f��q���J��{G��Ŕ��N��ܦ��|ڸ�[k,AL�`�18:.n�3U��+�l[τu!��2`�(Y�ęf�1-�$A���K���A�L��v9�g��r�K���k$l�o'��{�A4��P��#��N�i�fR��=�D�nx�P�C���&�E��o�����"��/#T���	�,��g6̘����l��ǜo)��QZՂP7C9خ{���ǟ�6ʳ	�3��~�7R���G�FmG"�L�)¦l�]T'��Y��u�"�G�!˰B��u���y�HD��?�5Z����۾�d�"\���������m�c+��� �Y��kR7U䝢�� C,:Z0m9�c!Bھ:���+�Mޯ����	�I{��W�>V�Z��~�3`�	\Ny�ޚE糽����tG��������w��h��b�c�-col�ޞsv���M3����$�����&��Sk�ӟO���]u���$%>��L�\e�y���� �[55$t0j�	/ "������+���R�O���������]�q��"�b�R|m���#Q,���ӒWw���zki�������geHƽ�@�����T��s����YuE��đ�����	�iKv�6�N�E�y��9�O��Ig�JӾ�*V�5CU������[����
�"�!�?M�&&�sg"*�g:��k,$����RYl�91c��ʇ��2aܿT>����a�1�ɼ�#�v���ȳ�_��w���$���vR����a;����}h��?�Ȯ�9�ɱ$����N{�"iA߶�;ϐ�;ka��8ż�y�4�:O�	F��9B��h*�ku~wX�4���j��k�$6J�
�+����^柧ַ@��;�F"�D��ȸ�XA�.������!BC������Wf,g������a Z����Ӓ�8�b	�hc����(%���1s�,�"K�������=ũ��������bU���=d�R����JSǯ�Ҷ�*�%Yú5����[����F	�L;���_�t��p
*�jӲvB�`#>?[�׼ʚo���Q\�� >���s��Oc3��x!M�p�E����A"�k�����@A'�@9�[(��h�2.?5'dcw�>e"
H6�V.��1�� Ff-8.k�q�y��	Q��t~��9���e���jX|b_M'쩀�����L�u��{�i<q����Kc6�:��h:ʆ����#Ӿ�2���F����%3T�x��È����,<<���e��d�`I	����1KKK�C\���a2P�b�ߡ�^�,ŒYcኹ>Sُ�u&�Hzn�f�<�b��OR�7=RX_6���O��Y����9~=r�6O1߈Ane]��g ����/aL�X�ec@�M?B�U�P���VL��:�����IK҉*!�}�W�/[ (o���0���f��sl����4�5&vAZ��L���Вɋ�'Y�؎��G�^heķ�[�؊�TT���4�0�o��F���0ky����B�'֥N�U�U㇧�T6k������*n
�����xgbSA?�%(j�v_�Ì�����D(f+�--}f�������@�8�N2���W'	M�;͊��O�LT� (��B@�'���$�
�J�j�.=p��Ҳ'@�.���i�5\sHQ��g��L���K�ᨘ�p�W'���3�f��#�Y2�k��g��k�I�Q���d'8�3eMWC��WF���L5Ϯ��f�;����]�'������N%�X��r�s���� ��iX��E��y�R�L��"J���e/��I\d"�{�$7����/�oF��r�b꺌_��\��̰�^L:�Q_J&4#�_�Id%���a��>?A��*_�AK1�Y���y���x���m�÷t	d��i��JL�ʳ(���5�V2�z8�G�f]�fn	$��^4hM���
k[5�*X	>��X9`O/u$&&zl�K����ms�K��P0m�}�z�cH�sz�����Y�f�[;e�b��ZV�������Lo͙iܰhĚ�'_���O�v����X6�d!���k���$i�Z�I��߶+rɢ��V��mC{��y"�B��=X88��c�*���Mf�hhi��P$?�`��H��_��_�,�;4�z��� �w5v�����t�E��4�;�ȃ�m2٥���4T"��Wkä���^��Yx���E�@P���[N�Bފ�[c".�L�/��t_����x_p�3�vȉu�D���i��������n`1_��%�;[ >%ϸd
xhd+F�,��V{�mi���Xj	�m:)��_[`fF�!'�c=s0<g;�}j�6�\�\A~>���i�k	P�MY��K�(If�Өkjtt�$�W����(������12��N�l�������C������W�ԠQdd���~�ӓϾ���a���B˜����:�{����]R��D�}j�.��^̪�e���QY��J��,�B�������]��x;�Iy �m����Ef9/�iK���ㄏ֟P`G�4����>��\cm�X�=�ļ�k���),^©k��6��5�S��Cϝ�`!Z�]"Ck��A�}"�gıU�9�Z3�Xu�J<}�"�jb�J�����N~�d�2t�r/���y9j�2t"f������~u�N���&L'"�5@��ѻc(^�¢,���y�Oh]�p$"�%�ܟ�V����._��3r~��ԭ�"t4I��c� *Q�aíf�D�vPnE���3;��^����2H���G��{��%�r�,(A��ЕzmX���⣕�Da�PTj�A���YQ�4�uw��/���F��Ȕ�sS 8sxh�֊ə3l�"Y(bfF�Y�U���Z� C�����}�O�5]������^�18m|7���$ۍ���L� *�*#���?���?���$?	��2P.1[�f~B���Q8�>�&����Q�pnʨ�T�~��}>F��j�N|`��#}B���OGO��?�� rlH6���p9�ՃTRf�
=�1��7�������9���M�{:�ȴ�ه�֮�x���ZMB��/�=�-���T���~��y�"��؈6��"qDKR�f��Vop�if�g*���ċ�|�}uqq�9�m���g"D�
� 9�RZ]���b.i�l`d�Fytz�nC����ϟ?�zRN���
xr{�H+ha0�?��@vm'�(��;� G�?���W�ܬ�Ǚ��z���N�Z�t�Q��=�-r^֒�.nn�������6��E�B�.Y_�ev�����D�����IĦ��g*�*��j��i�
�-f�R�xb���c�QE}q�ǟ�t��]���{v�r�)X��u�p���b���^DLj�T���ǲ�D.m��:m�ްm2G*bX�P7�7}x�BL�$2G�l�J��+�+X=6��7���b�C�l<P̡�|/���=�G�D~]�ۺf�m[�W�3��G����@��ʓ�H�_���=;;K$5�OS�ޭ�as�}��䜽��#�t!����b�j6[NBk�գ��֠ٶ����TH�f��o����k���p��,v�bȨey���L�_+��mΠN:�%W��/{�r��}ٶ9I����	>t�,��[��U]�{x>�	�!�y�P��aEix���qx�������K�oT����S�١�6:Igehڀt3̷��n2^�J;!�*�,����z�8����l]��]�8���hmo��8t�{J )M�/�l�`��w����$�T
��_/@�i�!�]��OQi�8qO���@7��8Hf�9��}�;��Ђ%{�F(a���f�8��G�����VS�F�QTTԂ����@���C	뷴�%s6���@G�v����;J^Qls����z����[ƶ�=��V�g�^�k�P����Q�d�ٹ9 ,\�Թ����;ϯ��V�*Ls/��ۦ5oY����ԩz�j�<!�(Q���2ͷ.�F>.(��$A�`)
ц�z n}A3ں��%����qg��eΧ)�i���8c���̠^�i����pH|��3��3�t���S���BD7ѷ��z��4D���-�h��n��[���-�~7���l�����y�K��{�tE2R�t��p�}oO5LD%	��6���u;�eX�0�)��~����f��-�7������>�穖������������Ε@D[��e��o޾��
�M�����3���]N���
���(���M�g�[�~_	��` '�Q_o�,M557�i�82���k�qZߪ��d�]�4,@]SG�:<ě��Tԅ��ڨ~���F;��� +◲�j�E�E�����P��c���f%���e$cD8��4i[�T/;�nW-Ƞ�7W�EM�׿|聯��=�?��Bvei���:H���z�W�$�ߺ�`z��*�2fU�ޡ��P�����W�B*����8�y�X�z���v�Bu�Bl���r���R��q͙���E�P�����*�m�@5��{㸦�uY�,��$Z�.��u���g��(�M�=p@�ts�8�՝lm5�C���n���d}>y�w?��"E����'���S�Q�cUַ����(n�kٿ�
�����L?X�S��k�IqA@cDJJJ
״�%�112acc��n8敗�����,�����Utt�Gv��[Z�R8��CE����;ѿ��N�����\��v�)kj���M�u
��O��iKUA�<�
�q�����@K�A����1���LW�^ 1��**G`�V�%A�y��6�,�3.�dr���ٚY�CQ`f���J�XT����#ϱ��یv��J�x�Xx𧗶/�I�3�~[ƭz��m�����Gd�������	�ڧ�Е��t��*�����k�yq�I<�F�(%��D==ڵvuA�RŬ*2"���uoh:����aC�|�İYn�{[�Q�QK/��bq����~+��c[k#B
�jl��Ēǀ�x��xU��z�0�-+�����Dttt��!���k.��� ���R1'KuN#�v�����b2|:�:��ߕ)��
ZZ��x��릂�V0/q�s�}���X�<��ff)��Yc"�ɷ�v�u(�Q��88yyy߆��)��>����=��]��Q��X����(`�L�`�>/=ݺm]#��L�o�喾��t��m�B�����ZR����[fַ��}��7�S����G�W�nJ�����e�L�lʫ��]!/5=g;202u)��~�Q�Egs�g��̔┎�����fJی�p��A�3�JS��66���,�,P�F!�{JD쬅�xg�Ц<+��d���#f@B��i�%�����;�{��cR�x�MmYӃ!;��-�YnI˻�I���U�>Q&��Ce���H&�M��'A���Ywn3moqC�,��k"G���ݽ��h(ф�9��M?f�/�7��%@a��fcd.�J��U��DBvDuu3g��,����M[�ې+�W�����Pi��2�CFLe� ms\u]�5�lO�.j����K������܎��M6	7}�����7��WXG8����#�����J�_զ����?3-�2K]�K
i,�U,M��~�>�C����ٔ���Cvna>��!W;���K��#%��\�ԾH����^�ϖX�t�}}A��~q�E@)�T�E�Ё:�3;?g��E�����W6N��,U} �������,ʆՓ���Ɛ�B�*p)3$�s��7��v�C�ֿw�{zq�zܐ��UVM�����O���(M,9�N������w,��%P�E�C�i� ����(��lQ�b6����hjm�d��L�3|ІQ740�[=��	#۽�2t8�,�������`3mF\���$�ϟ#mj:S���ne�cF���q�M�0���o�Vv
O9��u9���.P9å���<*d��0�m+(A^38�.�Ҹ�(�F�ˤ"�����ͯa~�U,+��@5����~=M�i��'�v�������sT�M�:xʱ�V�rlEl3��A����]��[׷A�j�3����>]=��|omg�����x���|-d��Ys�����U���Z��n��gg�M�\��)�"�G���_����<�pʣS�9��r�bs�Nƙ7���!�7N�X�x0�}������2J�؝���V��)ur�F� � �B�(��"�|�@uĭf!j�w\٥9o;��m��E�!��y_J��Ϭ���ue�6A��'"�k�I��*���/!kGR2�k�\J��hW����c��\�w�D{j�� � �)}��Jԣ]��!�gK�s�=�O��΄����S�%%ZL�j]�ڪ@�?G$۬�@N �����H�P���7��>#����n��~>��9�&�o��X{�	��F��0.� sc�>j(dM�r�4`�I.�E�|����RuV�� ?��x@��b���f,����-u&�w�z�<���|ASGqv�l1�$i]u��	�r���s�쎼��bQ�$�V�|����#�8�D�¨CQ����Ixz hQma6 �D��c��[�3���>>�:���\\�j7JЯ����[��������Q�����;^R�O����3��4�d�s�E^m����/�H����.�i����M�"��Q�g�E�%��g��U���{E�&Xٚ/�^���^� ��2�苷�����$`�xkn!*"�2�$�fR�D���m7�p���_����7��N��JK����c��$�/��'�u)�R���,T��G�G�7̭�Og/C��qL^@p�w���QP�l{�v"B�\��?�^8�?�����!5O�G�L=\�"�Ϫ��j���Q*[1�.a�h Pm�0��pS|I�C������F�Os%{��W��Ts,�U��o�W�G5L
f�	[;���d�ڹ}�nlygk�%{���g�T�8���]5�(�x7��x�� �
� �U�4q�щ��nOH��w���|�KwL �u"��O�ͥ	��9�)���O�Y�E���:��1�vZ䡗�۝��*�-�a�+�-f�BN��,l ���I^�d����7
cX�v������+Kv	H�Ui��T�CXdG�� ~�����=�uj`S��>;���:mN�0���'8��彂���_rQ������r`�R-Y�Y�M���+���,a��������St�+�X76���I)R��L׳�.--�n�oI��	ڒi�gwuA���+�)N���$I�wÏz��tb,3���L}eT�M�6R���t	H7Hw�t�tIwwHwKK7H#!"�]�%��\�ϻַ��C�ff�}�̜3Hp��+��f%�?������I�*51����(3�$GAiP�R�U�X��2��KO	�<ė3o���Dx������>���67B\�8����p=��p!�Pt�� =/<Mj�Y���!U H+mݞ�hq��	l�Pa��d��p��)�&�B.\�'"k�kO�a�n��WS=?R�\/�}fuK|�!3~r�����[���F�0�ߟ�W�פ�z53R�Y�}q����	ج�`��QKw����#0F0 9�jl���N$�0w����^ZN�633r�=W��GD�߿�%&>�.�Z���aS�t\x�p��-�T�a��'�H�	�^{���tw���+ǆ�l����J"�|�F8Xs!�C��v��s��/鑉����V��r�����+��^|WÄuY�Xq��wi�=;�c��}V�y2�%Ȃ8c���Y4D&
��^ �d�ΙC�+�����×VL�Ì?�SБ�~����K�>>����4�PbحƮM�
_,�����%N;��x�<?��}o@�^/��b�s_�˼t���;pGb5@��O>	��t��N��$q�Hi�u���|;G���D�E�����O5'�k,�-I�Zc�b9��DX��2�PQS1a(���*�ſ\����U���w�,X�\S�ڨM�Ĕ���_lɦ��|R�#��L��L8�	��c���L�$=g�q�e����C/
'	#c�9�iG��]���}�=	2Z��JN���˷�Gn�Y�-�)�n��|��q���>�I�{I*Z �+$�k���}݃��c�lL[���<⳩����R�Ʊ�4C�ɽ�i��� s��}����<��v]	/���On�6��0�j��'����~�O�E��+D���=vu�����x���
B����D����rwA�0E���5��+<O#�ʬ��uDz���j ����!� �~�/�#�9�Ĵ��i��ܮug�r���ᚎ's�+�4NR�7��U� �܂v�M�-|^��p�lIwo^����P��7�js=I��5dVr�i���+��[��WC����s�!:��J{FrRL�<|�x��̓�}�o��9�*R+v�gK���e��&><+rQ!�J���TW�C�+���k�w�|��U�K E��S{����w�FCc�j�D^����/�e�/Rv΃@8�O~���.�o�ҜF�t��ЭecmƔ޻�2D�CO��i,	Fye5��b1�p3��q���OU��p����j�ٵQ3����)aa ��q��"�"�~��Ob�؆
V����[��㾬S%������g�HF��[K�?���P;R�_)�(G��'3�r�60��MOM�ڌ�)--M$ʑ�쮥������M`l��f&�Si���Rt(�m�v����>|t1ײ����M��8�l������/�hs�?}�ߞ��=Fzd8W�o�IZء|W9�[����#�4Z]��U��+���6�K�����7DoU���	��{6�e�kQ�`�_*���X8t�q�#L�,~y*L�k�Do�Y,2�UQ��V�v�8��f葤���@���i޳��R�"�Dq6}�Z��2��5Tm��ʕ��ʲЉV�،//����[uAtX5U3^31ӗn����O���0M+������ɚ�Y�{GGbJJJZ�I�˧�ֳ�;�c��%	{z�d��d�2�����x���3o��wփq�.�����-J���V�`Q)C����,�XZ$[B�ױ��ɕB{��$�d8���	"�Ԣ)�Vu�<b����͗Z�#���X���$	g0�M�1(6+yQ�,n��c�[�Q���H����[��,
>J7jԽ	a���g2��Y����&Nч;R�1��$I�U���/�6~�D�m�(Z<|*�=MV�|��*�7��_�o������� ��2w+�ީma<�K3!''糔k�!/o����4�RQ%��)ï��]�҄!�lxtɉ���s�B��*�(�xa�E�����@�l������tiV�6�YF�AO}H(lx��?k�cG�����&�rm:��ۦ�\(�.^(�|�?浏�d<M"�{P~���!k�RbJX�:gd�"_J9�";�`^1���i��Z[�2�r�[#"���}���X)JϑV�+~���ش�x��ɏ���6ǆ�pV�� 0�}��]Bh������~���8X�I90��d��Y�Z.����+�9��gcbR�z��مߙ�����UXb�Tk�C�3o׀eS�M�a�Vc�E�9e?ڪ������I�<Z"��U��DBG��l���IO��H@V��[A��]���\�u�&@x?;b(t=�m�-����8���U.��glȆȣsՈx���
A���Y�4���"�;�y#��q���$�0�>��=�i��#"��aۍF�K���0�&����v�[蛿F�"\\تm����H�E|�uև��^�QEG�k>�[�ۉ��j�ƽ/"� ��O�8d&�V���=�,���TmС�x7��7�A�x}o��܉�Et��+UH*��4���k�n4���P�_�Ǌ`D휉�\�� ��7{�Ұ��)P��Y����yt�����k�,��}Ԩ�o��ׂT.�62dƘC��1������e!�/}!=
S�;u8�Q��l��#��*�6��rD?}�$=�΅
Ô1R=o-��V|3\d�z�*M��6�-��u��ȦU�Y�ee>h�����J��|;�ye�{�sڞE�����Q��p��q;�r�S1jP.jR���y-�s�+H��O��pcE�So��~+��{�sC���y�mf3�'�h���\��DѨ�DJ�޹$�q�؂���eo �i��'���wT���A��v>P�^l�/};zy������>�K�z(�g�Б��TU���V���C��Mv����[��:(jiI�%��|�@$pG%۔��ϫh@)�2�z\��
�\�u!,v���4�eB�{�k�~"kX���\c1U��I��K�Jc��������<?��R��`��v-���3�)�����>ag�9��H���Yc!�L�`�㿽��e�:��
��,�.��ܣ�tu���:K�����G��B����G;v�3����;��X�\���8���QM4i�쭅3�
?C�o�������,�p�����Uӛ���t'8,h~`�/�>����"���:(�X�-��n�YJ��w��P٧r$P[�������ʶOǀ�m��k}���1/��No��w�PPȁn�<G�u�bJPP�}�l�G��F?��F�I�{���m4�m9oCl]����wdܩ��ۖ�7�,�T-�!@���^�Z+�OWk�)�ƁN'(WAGd�P�롕�I�By�aG�۞��6:Zh�z~8�,;˦�,��	g�#|K$$�	��暿{04����Y�`���/�Z�#f����|ji�F�Wj"��
4�_��
G����u�h�#QV��C��ϑ�ޟbj$�Y�z���2�)}(��`I�s���=��U2�����A�����_/b6�HR�9q���Y|qe�6@766�̈�&��G�`��g���
/�Đ�bH��{t�;���!&�����WL��������I�b���ڿ4Z�߫м�;������~Σ�y�ܵe��,��_/��Mx �8�-������f]Ã8� ���4��'�T�i�E~�����K.��3=N�➏�aC�a��=&��N��]�t���M����i7Ƚ~��ma��E����#n8����t���k ������Ϋ�@@�������8�n�!s��{Y}eee=����==�JF4�t�r6(5bK���Q�{j/O�y�a��p���]�(�K� R[R.|f�Ka�����o���HG�R)�t�I
�R�ɘ<6{>O93�35VÚ�����&���І�Qp%�i��*�<����������n331A�����#�E2��W������IPFPR��Ԥ�DDD�Ck����AwM�M�D����\����нJ������p-�f��л�Ewj`���b�F8��* >Ҷ��0x^L�~<���Z�0�_�^���+a���{�iY�.D���p4gl&��}u���*�xy��ð�Ӻ��j��ҿU�r�&�k=���'��^����5A�F��>�#�a ���q�����,T��7�eB,-}�NϜ!?��M��Eh��p�S;#[u�i��œ�G�2��B�����#A҅Ӗr�3 Wf�"U���kS{�y����Y��<=�G+䮕�z�8�m*�Sy��J]�P.���/Q)Q���Rm�2܂/��g�k��,��E�:#�3�������ݥ�࿿�>��C�+�8�n�^O\:��`B81���|&����w�fn�����?�{�vЯv��^��4�^��o�D-,�s��|\Q��@�M�d���Mx�p��GgΆ��@nP��WYY�2E2)ҍ7��m��PRPX�	��+>J'���;6x�AZgrDIʋ����gzj���`�+N��{�_����IK����<�t[Bt�ِf�8I�b�^Ƒ�[SG�+�ޭ0��J��Z���b=L�Z�㾻%����Si�+��Ր�����x�
wt����R��)���3�����>�U�b���Z��� [�^����ܐ�}��fdDKJڪ�e����+��NT�A��,#�vx�**��,j�"q�rU�W����7쩩t�W��s������X|N�*"�@|MH"<�ܕ��/�N%j�h���O���(���f~w���$3��y���vƅ�v���A2�VB�o��yu�-����A'N���L�9�uʒ����#3�����>}_�60��I�`�Z�M9b�6aIs�ԗ�,&����d�䤲�$ʩ[η�{��Ǐ�jC���}�Ȋ������}>nKDl��ow�΀St�
lN��}�J����;v��(�q����)�hM$��ᆕ6�Q
�"U�b�9�R�
���|�c�,)�"��>e�f�3�Ҝ� ��@���G����.}q�ZY]��wg��9yK���&�7~5�t�k�P�	R�׀����T���JhQ�>S#ss�8I�}&�|C6<C&��q�\��n���kY^"	�p�Sc����9�x%E/_��V�����(��N}�z��AqD��_x<v{]|
!A�a���n�����3!���e��I˧/;�M_����md,���^AX�����������uǠ�T���_�s�ƏXbJ��t�y���⸑��
�gD��'��ʡ�qu�ߔЫM�Oaذ��.�����E�o:|�Z������ٶ�#Ǚ0D9yw��WTD9��˄=8<�4m��ɞ+jhH**6�X�U�&))	�(�;Jb�lm��q�l��\�������?~�}j�I��lD
CٗpնȎ����ܰn~�瑒�j0�r�:ܸY��+�hlz�ę��=Em}ڟ;Y���q�;�]}C9�k���۰���i�n�xA7���&NfHI����#�{����&�AZAo�_f�r�|�hZ�Zb�Y+:;�!��LM��+�1s6j��LA�x������~S���E� Z���d�%k";���c�P&o���8ȇ����w�44���xBƩCBC�98(�چL�ml��&4)��~�{*�$��XX�e����.&�S-�J��W��ѥY��?n~68��чgA� �T�j`����9`���$~p.�ˤ!�~�\���PE���TA�T��k$�'�x��oa�Z9	^tE�Q	�K�j�B�ʖ�P�P���[����2�ٟ._������q ������:睲�T"���Nw�M�̋@�'�NYV4,���*���/m,	��5~�eM}S��,@	99�_f�5�]��q�֐�騱�M�gIR��F��~i����*a{v����VDLLl���P��.uQQQ׹�V$>�du��3�4��SM5UT�r�k�.�#�M,A��p��񀝩`�fyp-d���/O��kO"�LJg�Ġ �� �m$�`�k�0�C\�=T�b���mw"�[wtX�z��т��Hlza��<QoC^ �t�u��+a]���������;�w]ts|!�N� ;R,��3vɶ體������&m�w����2�w���w�#C������n��q�꼄~� 
Q �4`�rP���u�WRP9���DޭC���Ɇ���>p���\c�ig�P�5�X}b�Ohw3\0�3≇0���Zw��ܰ��-�҂\
Q�c�$�T��wEh]����A�L#�_�az�����9ٷ-IF8m��Ҝ3����9=��9�!/*/+K')X<	2 e���(��A�Ɨ�*�$���v�A���c�G��U�ې�룣#��AN�߉Z�5�čg�L@޺����8:�E����?����l{I����tP?�逌�ڳs^���0�|0c8�Ξ?3ۤA��М���uq�((��;%�g�\��w��g�2qٗ1b�����ؽ%me��y�Q�kތZ�f��o���y�B����_&���0�i�T������?ct,0�2i�ř`�֘�1.cT��^qN�֖�֨e�$�ktXң���.&d�J��:WuF[]���h`;UUߌ�ò"���
2����7f�PRQ��J���s�|�a�,%&P��W�9�q�а~ϫ+Y�ٟ|����h���ur����$h:X����3��}���K�ub�5-�X>�Wf����B|B��DL�wV�O��@�i۶X-E�W�/d��y�S�˦O~���d~e��]�<Ũ�^�����_,]w���113�l�Dl��<���y��sݶ�c����K\\B�c��������L�縉D���5G���5W.��+�HT^{M�g���5E�@���E��7��!���L�2�L�LX�Ν-
��Ť۟�O..�I���A�p�6� �Ԛ<c�Nɠ�}.�\ů��ɩ��\ŨWMMm���_��,bs V�ю6e����K��yњCV^��O�]o`c�H]�
���153si��e����� ��u��wjv����QbYY���	Z�ޮ�mw�ě������g��ݎq�)"]f�?�f�~���H��v����ؚ��9�gh���,aa�����q�t=q,��#��]�>$cTX��a��[A#��#����ō4��EQH�&�H�tttD��
���.�=�������*�#A@�4aѝ�֡Î��$�R�̫XnR����8dRK��9�@�XWWG�Nc�<S���
�ʥX ���2
�1�l������^@}�c433��?8�䞙�U��v%h���'r�"����m�p�Ӧ&�9$��?ʮ���z�w7���x����0�(�۳�m�S�j�E]�dV޽OuVXT�����7�pte�\�7��2���6/�Em�4W5��D2A,T��z-��{p��5��������g�ޞ���������Ç��S7FX!�ѝ���y&d�w qC^���.�Up�~V�DGGW�U�xx��.����1�}��j�.U+'���ՠ�+)k=X�ql����(yʰ������lO�{��^��I>rq		ȡ��T
��o��-_-�j�cH�]��\2��{����o c^i6:�%��)h����i��;�P&k*��r��+�/!Z<q0?я[�}`ïc���sP��/��������9��H�jii!���< %j����<�b=�����O@ۛ؁��fs�v���e�/~ ��b2�x�u%
���RD�sN~�3Ͼ
�򺩞6]f�\jX^QO0}��I4/x��Vغ*�-KTh���w� �6G���!����v��� T� �/�����k�,y�.�)��6}�L�P�?��É����.B�]��?�}z��]A�Ѕ���������O���O�8��:��A�y��]��HY�hV�E�a'nx���҃�֫�8�7&&&..���i:�?�+LL4C�G~k���x��V���j�?n��Y�a6T�ji�_��,jӞu@�ͅ��� �D��_+����*\��\qWγ��VC�����s�i[�J�}:�D�=x�jO��YI��3{����~��n����٬�~f���FL���b�}�UC�&/bI|����YWE,����evZa��qq	�*l��0PC��ޛ��\^^:��󭶏��7��N7ڱ4��*aY��j����En�]|�Z
!%PL��!��j�X/��&I��Wv���$��r:hN�ƀ}�����^[��`lj�2I�T�Г������՜��jÛw����\��0�0�G�U*4����-[�d�����0|wق���<]�*״.�^���a-?~L��Y��pM�^ |�;�׫�}�_��5�$�暡�W!ezU8��.�3��ɦ�~�Z��9���������q>u#�1!a�������㇩�r�_(�z�{C��Q����$5t��� �ٹʶ�I��*���!�?r�}��t�;D���*�'�ݸ��I���G�L�K�7,��[������͏'��]�k�e�(�.dd�o�C6+N�p��u��q�=�0!73|G�7#(=����v~���[ع$�BB�BM�}S�̑�&@-�y����_ �m5e���w�h<�����xi��뉽�iS�8I�<��}��/@\sdl������ՙt����,�������g����f@ �@"��1(�n���s�6���d��	�?8k�<�q
�x�gɄ9����P"׏�<˨��!�8�u���¼F��6�b��h�7.m��s�yUUh�$)#�Q" )�&�I�^�������rgѿZ���CG���ʔWT}S��J��5<<<��h�����F����??�z���Q�� ����t�Dž�d��9��gw ��B5�$>Z������7D���	eߛ�M3�'῰�FG~��~OE��z�fIw,
�B�s�᪈�QǣT>�� ���t�҆���\��eqROahi�������+k.��؞� �?[|#*&ƅ�%����+cݼujjjukԢY�bMM�[xy}}b/~b�8^��U��Se�A��>�c�6=�j&3{��%|Lh+�V�M����&���7�D�5�C��(���jɟ8�8��:���<��)�\��h=L:yN�]r��.�3:�O������喰�5X�=���v2�k�$)��'�uf�F�䩎[>8�B���J�2F������i�s���<�kYR�d�^&�F���C�`p�F�Pd���K���~���l����x�+!Ղj�_�
�In�o�'�~+��:;��_m������P�����j�m�?ɐZ��]��)}�g�N#緢�S������w��WvE��� �*u��{>lQ�(�PH�������9�X7�@���ud����⸗�|w[�:��}w��v�:\�l<E�f���T�����v��R���(�dS7^��2$����9f�Cc�^�륺�C �R�قKE>��WiUl�,���p��|�Ž�\Vy�䄲���aU�E�m5hs�V8�3o����`�����NE�b�-��xuN'6���N���^��|��'�k[�F#H`�n���h�8k������X���B��+�w����9�s�Z:co��}������<�Z�7iG��'׽fuG�����7c��A����Ӷ�Lf'���<P_9>B4[��hןg��޶��6��դ	^���\� �O.D���"��xbs�|����q������؟�������pT�ٵtOk��
��|�����)��0�@�R�,�RK��\��Mi�5nV��C&��nOj,�[8�#JhN�_��Ź'�����aJU~�\��L^��X�<���*k�~�z#�ċ
�_0��;�����.FTLt��Z[�F�~����Y����G��]i���Ǌ�C;am}�]4!�]���A�l.X!%C�}�ȗ��r�+�������aO$A��zxil��|�'�pQ���aa�����;��^�ꍋ�֯���Cs�D2"~�?�l��Q�4��jĬ7�@blu56�68�zaϥ�lS�i�n�i����S�_�.���9���ʥA�-^rn��c�=����y�2�]y�*�"��⍜3:@�\,��?��@b`o����i�~B��|��N�{��S�M�?�>���(�s��c��˵nUd@�7OG�0;����o�̆���l���)�d�X��`�� $��a������뷊JC�#c��dI�ӆ*o�������k�"�O��1���E���|pt֚���>?�W0H��s�~S><���
z�r��*pW����BQB!�Y�AvT�w�∟x1�@	xF��
�S�P����3,R��ˠ��gr;_4���}尰L6���[F{]�йP�O��de���J
����jΘ/��|݉Z�?�JR����j���P�S���;�� ��v��s���AG��|��yj��5v�Z4?A+^�ɕ%߬S��. �+g����z�+��g�jq�D��߅
��f�3 �3��{���-��h�l���"#�����B*�q5P-Eئ���6����S�+��`�>�V�*/�]\_��6�猺~[\�9_��.O�E��՘XRh��D�D���n��-~����aTù������ w��F�&I�і�)��g������a��@/�@dR���v�p���~k�v7�i��aȍ�2^S���/�	��������}$'
l��޹/�ν �{�� ք����c"��n��N�;�D&C�p��n��D�����+>�ZEEI����_X����k��zOe�q�<p���Ԡ7L�A���ǘ�eZh�fF���9��'��������xLp�I�g�-�ѻ�5��6�h>�a����/�r����v�A�'���y�V�ݽ]�K�y�hV䞶�<'�Զb�����,��� ���E�aGI���82~a�dSY�t����_Fw�=�[��|����:�7�����w�>�N�G���h��/ݠu��֪�57�& L�m��覞��4��Pbܲ�ƒ�Er�����pP�lGE�w�o'r��9jQ	uދ�����E�/�Ĳ�V'׌%7ۍ������CC�)�����gϩы�m9���$�p��vG��ͣO&�t(�8�w�ʴ0�t�L�0��U/�b~ǉ.�|�KQ�A}�#�:ō���#��R��^��I����d3�I����B�XY'Ϯ����y8��'�t4�~�F*�y���|����_���ی���d�,�k5l���QM]ئD�6���e6�h��=!��:�;�����G=]kP�J��M<�o��z���fe��N7w����l�n��5ˆ��;��Z��Ԣ󉣬�>��� U[�?�����"H��z��ԍ���QQ�y�|޿�:�:�o)P����r���6��q	�mҜ�>W�"͑%yH��z���ɔ��D��/.�H�#X��ıd߬�T.D>�\��&ag��qij+�\�g�:�q"T��߱�N(z���N>��E/z�k{M9u��!������i�)ˆ�*�/���((Η:��4oD�ʇw��]�ږm���P���©�� ��G�ƺz��f���!�;6���E�1�~�.4������}'���g�Ы�����Τ�~��P�S�F�@�����]��e�;����e�R�D�J0HϺs�����g��lj�~��^fT3��n[�A�1�)���Q���S_�M��H{��Ŷ�U�~������D	4`2w~�djc�bee��b�^Li͞+��RF>QV^~#N��;�\���YYHH(7���_֖��ۗ�����w�7����.��ţ�kF��3��~׾r�Ȳq�7���}	9~[�-_�=Ij���aj�i5~�~=������Mv�tJ�^��2�6iѝ�x�F���6���(� �xu��R�
��%�-��p
).�."�è��ܞ��C#G��z�hˆ�d�����"[���>��y3���H����-��k9�ׄ�=��Cu� �q}��IS8,�����\��F#��@�s!�~�������OˁY�� L*��ϓ��)gGv�����m�x@)6n�60`�EI�Bm�ܤ(�����'�4�iK�g�E�,y�j]��?�c���.�&�����.=�-�z�����[�Y����T"����@�m����XGv�Ek���� �O�w�c?K��i�.�����z�����t8����2�1vv2����y�o.q�a�
]�W�b))�:�Kˮ�(B�D����a��tg�Fw↷���?���B�Pl<��V0���ufN�]�BU���E@=����3Ӯ����]�f{��&�k�vӆc���&ʢ��i=j,{�c�\^F/|��[!]M�E�&Ȕ+H�{Q����:E�;�r�<�ɷd�콕$���d�s��Y����]�3�Vxj�j�?��*���3n��>���XO�����n���#�P�Ypy^ѱ�Yi���ͯ9��R#�h�ڪ�Z�9�JT��**便]�@�6���k[�����O�.q��9q��s�S�h��9���;��T (�5��ԓ!����nx�<�P�e\uUը��\���
��֘�$�oU"�ֹ� �6'tg�[	���V��R[_̔'V���]JQbI϶Ĝ����OM��1�:H/TF��,��Eh�N���}�p>��p{N��Y�w�l�z�up��V�X]�g�2��0� ���z��Se��ඣd��	!1s�G�X��X�&��v�I�㥖��ӷy���PD�;�Y{���S���S��>�9����7�������9"���;+���Ř��@zs���H�cW��H��~�~(Fx|F*�Z�W6O ��N�h灕qr�$���4!b��[����?��������
SN�O���d�
f�������p��&-tZ�J�IvON����w2�&6a	7g��h_�GҶ31��L-�!Z&��4�xE��t�`ۻ���rF�ʻm���Lp�0>~�q�f�>i{.1}K^@��Gd�I���V��$c����E\��&��n�9�?���ko��O~�ԺcG�z露y�V�(�,���[/"�r�d��0��{)�����s��lҋ���	)��@���Ϻ��˳��qqqɣir���'? �VƑ��/�X(}��MC�eޚP�*�9��='<�)��ۤ<P��BI�-��3�q��"��o	��mtef�A^�8�Q��<Ee�+��Ƀ��G�^��w)�7�е7VC�`'P�Sq�/�޻��0<�Jc��Ҳ�=c�1�S��8l�7�3��,;�S�y4?P���Yˀ�A��.5�ǌ�ȁ8-[��q��23;���N�)1� �JY�/73��1�����TgW7o�K��7v���5'kkt��l��k�/��^&��rq���?ʪgdv:��W2)�$|�>�3p�"���t~o�-����ccƎ���|��-K73�µ*B�cـ�ˤ��/�֮���/'
�����	9km�V	�<�j�ڵ{]���?|������#C�TE�B����'//*��,ו������v:#C����aM�|�+W��W�<�ki#/{�����F;�?^�^��۷0}`�o.����W-Y�ˈ	O���܊�ea�^�Ғ΢�������<o�_�{����B�FW���NKLVA��𗕯vSL\�����It�?�0�[Z����8�$a]Wܩ�[v��z���໴��q��������p�C]4#��|����o4_����[�濂4_��o(�X�0'd��wk�d��G�����L�,E[�p�^� �ggg�#p�m��F�j�*��PA�yf_,��xc~���L����ǝ<�|Z�v���R�_J�/,�@���As]�愴��&k�3����C�ԍ5r6}c��5�@z�(2�p�#8e�?|J��x8�7�r�'utX��V�RW_�hE��&JJ*n��<�
�V"1kr������a��Wl'�W����l�W�i�^�`�;�9������>#���fRUUff���NNΚ�ߗf0iyH#�]<�Q-�f��b!�������?*�UG�E.`���YM٢L�NQ�OY���z����:�$ ��/��a]�"s'��+N� eP>�R���f��;q�dp�:iTL��I&4��('����o-�   �]N�׀�4���Y$<U_u�V�Zr��"̚��-���	~5�s���ᐂ��d�?�Q&t/,�I*��4i/fD�w�6�n��_z0��D�|�� ��0����v�-�t��t�9������w��U��a���?�YITd!���g��3�o���jq&_��S�Jv��h��������l�ZIN	d�p���<��*�����jv;3Z4�Я7�y&1�}<<D����6	8��;������[t�zrRG��Ч ʝ�[Z�?d���O�:8"���޹>�Y�vܳ�k>�\Y�ffㅍ��q�f�قlw�����Z���L�Mq�4��w@.`���	�������c�|6OF`_w��๵D8���ĸ��w[y�*�n�n�ݬ��9bf[�*7���;8�[mX�=��n��G�7�.���	'�J��N����R6M�s�)Xx`��~_�0bBC!��h�!��,6��|=n�0Gt>�"�1}���t�ϳ���rf��cd�� ׉����������S?�ؑ! ��\�=Wo��=c�`�Ě���"~��3Sl�Wf����2U�Ԍ�Ċ���0!���ܠ����j�5�"��v;E�T�Ca1B �f2�c]�n�v�s��S��Z�EU���\ ���KAW�`��B'�x�п�G�]���o�F�}���y�JYd�� �5)w3쌓;(˂����1��Y��0R�H ������@*�1�wD��L-
/x���A8����X������	q����RmҦn��T�5v�Ze�7�X�����y�53X!Aܮ�1��+� O��J)�_RGI�}�{$��E2�_��$
���`����y&�!~�"q�~�&��d�4��r��@��	��U�m˄��lr_?ZX[[����"�Y^^���3P(�R��j���a�>Ɔb��|����E�����4_���Eޗ���W�Ӽ��5; ��=�1��C��;p O �
���9\Z�X����V�
����O�w�����N��������`6?���3�!Պ��{x<@��EԤ�w#��s�y�"���9�M��*4a�!��jǙ�|�^��������;@��V�ȗ��&�?���SY����i���9---}�w�0B蕈�Mv˯���TU�	6rt|�Y�N�m��97�7Gϳ/�t������"^�4z�#vz�ר�_����]�9��6	O�����~i�o^�j�?�������a	�H�ݤ��n3ĕ�)B��2����^�B���ןD�0�s�/.�{�C��1��>���tb��xe�ɫA��
J�	�ѓ��EbW�\�����pDH',-�	��V��t�{�@����sa��6��Z(��z� ��j�ϴ¾��K�]�a��燪���.��^���1�~�DEdw���F8$�8Qk�:r����VQIIo�UT\n}f��,�����eJ������jsD���VA��5�<�� %�����wӱ����� \�bb����v�F)E�*���AFF֘A�Y׫R[w��xx9�[?��?إ�����̵r���ۖ�Y���x�:��̓�1��X��sF?���[SF�D�<M�i�ǄL� �������-�}I���L��}A"A����2q	�����ԙ��ӦG�{� %}a]ږ����zŝ`�/��
��x0@�ᤘ{S+�b�������>$���KQ/]���r��!|�c�@G~I_.5�F��H�)���rx߼в!�c$���{Þ����i�� �$���|	G���_M�ʁ�(�1+v7�;��S����<P��W��LA���xa����7�O��Ϧ�w:���zE�2�ڽnY��	�I� e�1$�\��hd�L�ny���*��#ʣu���#���Xu�`�f}s��|�b��s�Pi��8���l��,_��<��v<��'��v��]m$so���_���nyƐ�-PK�g�����C�/�����v�tt�����/<� v�HȐ�ü�N�T��\^:�	����9A�*"[k������ Y���}i�j�ʂ:,��bwc8{u^��F5a�XC����ў�:�VY��Ju���m�˨��[5Rs�f�םoz�	۷T0�RA�*���7�P{ſg�d�1�;�#g�A�� u@e���}c(&�E�t��ɉ;Z���JAPC
K4����kY������i�-"@U�.�4�} VÉ&4��FY�';��;�yzu����5o���U����G��4�/h����Ha3.T��`x�����޹l)��NV��"A6�?	�Z/e��Ԥ-�Z�k�A��7s�:o�=o��.�2��a2pTA�*Z�(<P3�$PU��߉���O6{\�<�	�Y�!���$Upk+�3g'���)n��6�%��&�L��n�#��e	{&��j(]�\�;�������K��!!���@�����<f���,qK����l&u����"Ŷ�o�<��}קI�xڡf!@�_�u=��زv�V��k�k�LC�v�C/�� �;��g�I����>��}�f���紪w���a��ꕌv�E��J}�U$;5�����U�����b������}���[�Xb�kc$d�q��A�jt�qR���*Qc�������Q�I"n�:��w�8 ��"s6��iK&�۳i A����UT�؁�ʥFU�
T�"��Z�^�:!%��2��IDUռ2�W��mO��Wӕ�C����5hbFB�a�%	I�ʾɖ$�-$
/Ë��-B�RT��McP����ʾ�R2D�%�sg��s���s��{��{����|�{�PfW��Z��"t����ְ� �Y{qO2��rO�N����;��%;�}�J�j��v�1���4,�D�+�����6��@&��ߌ0��zv#Ɍ����,N|�~#����p
��B�T�ͮ�!��%�r�}��&���Ķ&7��Y;"-�kGdF���}�2m�ɺq�'J�Y�����ɂwz��*�(m��K�>;*��?�����{�/�*OR��������ͅ-�]Z	���0W�Z辇��SQ�HA/��>���C���%�b�(�/���A�L]���C���:x����R��H/�Y<$HF"�W"���Y���D�3%�AP��^�J���b��d�5�Gw@SL�L	>�%�5�G|ڲ��+qUn�ާ�>.�hG�S�F!9�;���sA��3�hN�F�&�|����w00�^	���lf�lV��`(�,U��wx�s�{�>3�l)\��Kq>.d��v��=F�%�4y�ƾ�ǜǋ�փIz��퐀����=�<_מu���8��Y���������q�y���uʆ����o�Z�]�*�f�+ET��r��Ņ�@�<;+[�2��X����ؙ?W���l��!�,����]W��L��h�p>9[OcO�������:N���Xf�t�_��	�5��;I:G�[
�V��ע�G}j_����p�3 � '�h�{�^��{)Z�o�OҒ��+ �v2�D5~S'����-�ࡨ_�bV��[)4�=L6�\�g�
p�s=S�h�cc��uF/��f�;^:�#����F-P�Hӏ����Մ��&���8,�����4Ӻh�$JVI�n���h����`<��O��%XǙ��# �~�7fLt�n��Y�]�,�9�F9�v���Ո^�J��x ����}-|j�ʣr������ِe �/���3y�����f�s%UG6R�-#��3����ᡅU잸�\D�ջ%�(�D@��C"p+>)���yB�B �5�|�K� `�s ���\�N�-P0��Y�@Bv�V�d���	l���Ӹ��K`kY�>r�i�bw�FxQ�N�n���1��hS���L3Iy�_��y.��.��f���%��ϭf��Wfn�׉��9XѦ�^F���_s2�Y����-d{i��P3����o�i��f����~q� ��5҃Ěl���]!g���I�>�*�d{��R�*�%�E�_�H1f��È�5����&ä~�?���t�5QׄS��
/���qz�H�ޚi�kV�
���Mj�<c���B�W~�
�c���}	��y,d������	䀥'��̇�E�b�r�w�p+���{5�tHD��3�f�+�Q�	����R�=x'9w��y��ug��q�z"yj��HwL�a��.�Z�`�T�i#�ϝ(�"���͑�Arӟ�h�v�@��Q��U�+	$�ٮ���X�F��M�ע_巿x��Xr�Y�>�7�H�e��[�]^9s�Ӟ��K�����U�7ل��1�V�oGu'��r��ڛ��Eq�oμ�V��J��;�o��װ�?��!����[88�v��*�d\�4హ���������PeʧAn�C����ł%㛶�J��@�l�a��!m����b��_:�G�Wl�=�@��
O���A;}=�X~*��"������o��e��Ǔ�vl�����6$y�m\Q��Q�QS��J TMm�tDLC�Shj�sږ���7�E�F�.�J$,
 �<�R�F���4Dʘ�؎Q͝�,q"30��[���Ⱥ� ����s�$D�	���,�o|�nd�����4��l�6�E7Dq}��%����!���D�Hm���jSi8�`[r�]Ƣm��k�����5�揦�"��y~T�2�j2��Bt�������ݧLQ�>vӓ�ᠫ���A�z=��
 �`��U#us�!FC�{s��MqBbbd�n)8 ��|�=��_�S��v���-q�)Y�p �(=5�Sny�6�� p!��u�L��њQ�	^���v�`�f讀�j}^��[�,����k^c�` S	|	ޡ��,��>��WCo��g�s�1�8�V�xW �A�x���P�<���֗=_=���D�c|��V�j�X����@���,���ߵ�4�~7�kemʚPz���f�X�T���מ��`m��>������g5�3�0�*��p]���1VRH�6���VOT�5�7sTTeJ�����T��;U-'���:�4��ɭ�Q3��뚤N�,Ve:#����DT�~l|������)5˿�iV�G}�������{��ۛu�ʀ�_9�9a�Fh�'�xQ��ҟ��sG��a%�?J������vH;�m�հ%�
x�};� 쫃�����h_
������P-�0�+�c�Sc����DE�'��n5�i�A�0��|���Z�k�'?���+i��}G�.�0��l��5���[�a�&��r���h���튓L<����}��A���bo�ދ���W��������SZ\g{��d�*��*=��!�.V�'d� �r���@w��ѐ��l�%:+�a�9�y.[u�Nu�f�Lq���H=3���O�k9�P���e"���5��� �A��4�����8t�"���������P��?��'�;S:L�U 2��U�I Q�G�u�SJ���6��?�x��vQ���]lv#�J.=ATl�5�q��c�_.�	4�5�Y��l'2с�cW-RvQyeW�7�z���yڍp�ʾ�pᎍG1�A2��7�k�h���#MO�7-��9�0��B�������k�����;��;dk�2x)���T���� �8�"�-�b�����Ǆ8��p*�w��.:���?C�G>�t&�V��ޓy�@b�6��Q�,/���_a/
�Fʟ4:.u/='�0|��'#�0>4w9	�`%%CN�Ƽ~��aC�+�%UP{%��0V��%$8�W�W�k]$M�8�`Mg%>��ѧG�>��}1�p�;v���$pw4~��	l	泈 h�Y�m#�n�!��w{j�ҬU��8҈&�M�0=�HM��q��U;�Y���U��T�;�K�洜�!� �"00��z�[�AH꽈�a�iK~�0��c�1����u_堕LB��as��q�18��~��!񴡑�dv�-�1W_W}�J8ut��aa�����oAͷ���
�&y/?��6;(��#[ț�2�u�&��V�皣hj�.��n̡U<v�#Cw>�v-���\ꈳ�깞v��d�եĽzJpQ2螩@�N�̨��(�ɻ.�\&˯�������BI��.�� ��xh�xzP����T̄/��w����0�P�H�4�BF�\�������Fo�(x�AL�k�D(oF�J�1��l�!�� �8���]y���j�R�X�#�o¶��a�l��X|�zs>ξ�Xi��|$D�k�CP����ؒ��]�UJEȲ��]d����2��l��Y�J��=��Am���'>��8A+��&ov��_�>�Y{xٱ�l^|�$�������Q���������F��<�L}��[rXDIi�6|e\us�΂^��� ��	�3��>��ي�,<ǝIfZ�7�u|(��WI�ܶ���Uw���5o����Qa�Xv+v���K��:n�H�2��ݴ�U�yX)j����Gs��'R�Q;!�����9wv�	���'jψ�ԤNģ�/��{����H]��N�����Qo���Q�!:�X]˪~�A�x;����Y�d�3b4�bߓ�zx�:����N����ݞw�%�"Z��ڜ>��'2�p1g�Ca`37�2)6r��?PK   �a7YmS�;F� � /   images/45855a06-4846-4a51-b2b1-60b9838f281e.png��eP\m�&�2�'@���'������!��Np������w������TMͩ9��i���EyItTbTti)�2<9�2"��[$�����3̡����O�#������������)������'c{ۼ�:�0���b����v.0b�vn�N.�&��.��{,���$��=9�r��5Ɖ�~���U,��u������Y�|���ڳ�-��]{&�I��<XT���2_XT����!�H�k��H��)�E"�]{��P�$K�t�u��t�A�(�+=�x�j����� xK
�2~�&�w9�b�]JY,��nV��7E n4�<�:�1�я�������#������ؗ�3�\)�0SJ�6}�5 �!0���E��Vz��|�f��@��'��c�p:߷��T-�m�������ru��� �d���1j�+�>ŭ�3��!�/{�h�1B�0�m��R��L~�_B,�Ik�li]�(�:D"J(k$�6(O���x��HL��MZ4�4A�B`!t}�>YZ�Ț? �Q�@�Dy�Q�ۭRV�P��>)�Lgq薰�MA���@:�7��B���x Փ��a�Ӂ��Y�o�zϱ�(C�Z�潀�gB�P@�L?�h���׸3�î���w��������2���kr%���>��Z%T��ǂ6F�G����Q�!�����+c�#+�VC�	[�8�>'�C'�w�!�P�q��5�6�7�#�(iTšq������BE���/ Ȇ����uvB��a
��{��b�����@~��X�R�p�p#>�\�mR����P�4�J�G�w����� �ԥ�]�X�D�/�-]h�͌C�TR����.	1 �X�qw���޸��~��tC��Q�S�&Fۂ�1\��b-w�9Y�����Y*�U�e���C�N�X4Uj�Iړl�{���䩋�{�qSĊ]qm��K�Q.�2���r� B<�6
;{�55��G�� ��M�8(����@�:��ݎ�k���-�ŭ{=`>�.a�vtVk��\�_:��ȷ3�w�'���#RQ��`mlx�3
h�8���t�$#��4���=I2t#�S�t��Z&�
bK�@�L��
|���F�8<R�(�R������j	:���٪��Y-oߏ{ƍ&�]��%��Rţ�n������c�:~柔���΋��g=)/�v��j�0�\��	{$7�:0�H�c��lx'���o�MVH<�m�ɽH��5���?��S��p�m��y[�o�]����aa"��A�^t�S�.������w�v�,'W�E�`l���7c7z�G;����r� j7�m���X9�Z�1� �Q96����ϼ�ة�ߓH��t�����>��ml�s��Љ����&���|ɿG"6D;��̧Zl��yZNY/{����I&�}vcD�N&AM���D@�5p*�e����*����t�oJwz�)g�g/��_�b<��7�$>M~舙�6�0��I�\��;Q(�*�Z�M4��6��i����?�%�/�Hl�X@�L3�ɸdSO���<N6C5v̈́�޽���w�!�����T�uJ�0����-Ń�-��*L�c<"v�����W꾡���� [��G�e���Ň0�~���sw(������#�l퓔��\��z=[@ؙ��K7;�Fλ�#�0��������:B�����b����ο&L�)�D�,�1�}�"�C�~(i��M�Ƞ��Ιf��#)��0|��K��KBJK�)R��`���Z���?+B�-�����fI���0�1Wa���H�N�D2��	i�b�嘳�fKބUvK1q�������{�� �]Tj�<l߃R��-�|R�ИLBQ�eK�"��8n�]/go8�,�L�Z*F���ec*��"lP��>f�3�1�N��Rz`߫3�/ܝ��Sq0�4�=�F5�!��ĢP�}���f���%��x�*����)�?v�x[�����6���J�����|b�>�ّM��K�r���O�2/�	&�ߡ���I�������(�r+O�3��;�_]byU�dF��A�1 �r�����i�-_�Wn�F6��N6����E��\��l!��9�޼{AP�_����z&y2�_Z	V��7��	;�w���a
�[N���p�k=�d�%4�A�1Q�k��2�%I)"���g�͍z�%��fc#�ç�
�p;��!qȷ�|�5�w�҉9�=H�@������<��R�Zˈ��	ʔӎ��0U�'?���%g^]��y���P�*le6�R���I.O�����B�~����AIY*��I�۞T9�q���u��h�+z犯/��hI���w�[1gu�S=/.��[r����M�$	�V��J��5�TC�����q�*]^���Lv]����6�˱�h'�l�`/P����|�!;����6�$+�v?IFZ�܍�/���j&��x���b)��O�D��v�YWiY�>�+�2�b���:����/��wA���v�q��
�Bg����U8���I���_��`��~����y�|���k�P�֎��X�y���.��ږ*����wp�)��.<�� I.�l�D3�C̫���4�H�3�|
C�����l>���@��Ћ���7�Ǵ78�D+����B�[�j��0�����2q�U��.��ƕ�&��v���|��u�ʁ�J�Ձ��(�J'28;��Ȼ�ђ�]Fq�>}vD,�J�z�G�ᮅ�I>C��0��JW�E6aߩ�yK�e���>*7��W�l/R�B�{�;�G�r������_FutG�y�����p�DR��Ä�8�0��-S"�m+�M�io��w���H�8G�����<�������T/���@Q���,
�[�T��>K�ܯ=��1��L���[!�P4JS�c�ʔ��-��ia��E.��ߋ+�ȆiW�|��n��;�܄H�<�؜O�N��q-��GAQ0C���u��y�F6n��3_�Eo"�&�T��|"G�.xC?s�G�Gs9r�z�-�߭�z*qg�\(&�l~�pd-��ߺ��H�����x|��SH�uz�S�䊠����Zj���5�aL������2��G�`X?�s
�̛�Ž+To|�����:"�qf�كkH2|�"���*��D�����ը-b���QQI��[��l�Ae��	���� �!(����M�CUj�A�4�f}���
L^�f��tݱ�B�������䀁ǌ��a�Ʒ�\��u8��{��4��_�]���/�6�-DX������r~}yw�v�y�/��btěhFZ#17ф�nPo��/�=���mX�j'�n ��%k��OZ3��0W��/�癴�M�X�b�tvK�8q?� ��1:���Ɯ�`6��q�p�صN$��R�y���e����C��2�����'��ҕJ]֕�S7R�Mxo�|���md0�~^h�9�}2�e6t�5���L�Sö��Z�a�NI�SF�S��o�bt��`,T��o<Wұs���a�������RL)��SQf��dGz���\^�sf������6p�h�4y2���1��5D�p�6�hl�a�@9���y<����=14�� ������֋�N
y7z'���C��R�#Qxb2Țˮ�ב2�0F
���?�� d�o8�.c�M��׵%�Cey��a�8uU��z캛�ω��MlR9��r.&`�%�R����4|h4�jN��nLCc�I>O�;Ϗ��,����i�,E�C��31g��C�`��=D�!���Yg�M���j+�!��F֔���Thv��90f{�Μ+���s=C�����}B��9��wyT�K&y���a����8��-�ӥ�U�v!$%����2�4��!�,���%��-����k���W;՘fb+$��<�d3�8�ѠK 6�� �l�f�m�Л����%0ɢ݋7Ѥ�V�y��D�x�~���f�A!;�����
 PD�%�x\֝��&GV��9z�R�\S�H\��94>lz'�ec��޳���2A	W�r���)4Ht����X�j�����6\H����nH���6#�,��6��-u@uLj���8�$���f��f�b��o�$���Z�<1�����a�Ҹ���A?U*"�ݸm���6f��M_>�eE'�%���;l�~/�2�%�0P�I���)��ۼ�6�Dm��;�|�,�CD�-+���<��w^��񖁴��Z�f��``���(�3K�ߙ+b6F�Q2vB���_��]��P�f��X�����m��9j7�����m�6ǀ��4�ǉ��{(|�hUK7���eCl�6�^?F�[^��@���c���#���C6��R�#�V�N!��fȗ%�qO��������� ?��P�����bn����	K�2T���Qt� U'�-6��ÇQ��r[�D�3�n�>���q�?�]����t&��Gs̏�B@����=�����g������+Ġ������$�m�-:������_L�q!S��cݶ촛��>hPR��S���з��l�z��說r�j�\�k�Du�p���s�[� ���J�g�2y�t ԭ��{L�cޅ/����gFb_����ʟ�sy��<���N��[FI�R��|?���4wn���(`pccx(3O����B�@@z��P�ئ��7�Ɔj��z݀[%��]�*��yg+����+N����>+��kx���H����
O���e>\:��B)!Z�ߧ�;�x{{ >u��������M[
Bg7~�w��0X��LF0е��5�>̣�SB��7Y�����pJ�Q��ʵ�]��p���V�,1کx�^Mk��bz����m�O���,Zu�09I]��j����Yz7�[��4S"+s��I��W��4�S�UMܲx��n�`�YԐh9����+����<͛�=�C�]vL@%��B֩�w$?�jq0��{�
0"���y�����8�JCJ����4�\V%��
�Ɨ~��\yfpB�l����^�gN[�8J��}w��Ī�C,a�n#"r��O���4����\��7�v꿉��ゎ�r%y���q���Z����x�漀�*�_.B�b.�����NG{,_ �cq���2���%\��6U:+,cm>b?����(I����Dp[
�wk���</�o��n��(�1GW���8PQ����gxIB���7�tut/�S���6?=���t>�i)�.&Zƒ�G�������j/��"�2t��^�����qG_���#�HؔAkZ�^	���DO�(I�~ҽ��m��)?/����b(�����2����ц��&��1��%�4I>ϛ.������P�^�Іȭ��G�s��Cm�lO���n6�(�v½���tO��#?!�V�$3�'�����Ψ��줨�W����4��S�֙�Ht(Qs1m�I.T�0��P�������r阒B3D�^1�s���ح�x'k�מ|�yRt؊�P�\����/������ti7�fbΗ���m����U��/�v�\ԓk�a�\>�|����L�D̥��f���3K��F�W��'9%�{ysr�B+e`����������k��sL����G��4�P���߄\�������/�MWQ�,_��]=ɤ��`��HT����-r��˄��<��-��믯9��5|Rt�F7{������v����Ux e��8��g�'�tT�ݑ
L�t��{S��u��_��^Y*��_+RS�v,������N(Q�D/�N�@K�6��?��kG����4��A/!�w��K}n��ɊB��?�{��cr��W[/.9����ɓj����X z^I0��\a��G�:�f�
�C�����C��G9��H�4C��/��dZ�����w���NPM4�`R���S�,�o3��L1'���A.=��/��f؏�քoe�5׾�R�>���s0+a�_�q1h0ͳ��۠�� ���)�ȋ�5� ��t�t�2�󧩯�ErV���G�ME��խ~s�>:ϙ�g٦@��O��<>�K�+l�$����3���?F�[���+RV��t����4�縦�l��uU�nIMǄ��M���0���#�?Zz)}�,��"�eƗ�7�+%�#�S��"ym'{{ȷ����U�y���]P;�.����>$%�b/��L;��F���`��k�[%���)��S3��팛#��E�޽�f �3?A������ �-��. 2��4���'.nr/���������ƗH�/�{��m��"�Ac��K�,"$�IGƢ��0�Zz*I&���T�_)�Ǔ��_�x��=I#��C0�v+`��]v��G�bA��Aٽ:(Hi<OH�ހ�w�FN���O��AR}Ex"9��$��_�y��Ov���Ҽ�C�_)���_���{�N�Pk5ؒ%�A�����������s,,���4���c��$�H	9�t�xn��w�|�k1\�*o�t�)�y��1�hd���=�mlQ���!FG�Z�R�~�����^NaI�ln-��	���_�_����c%e~� Y$�Ъ��L�������ޡ���Y(�lz�%t_�6�H<��2B��}�]Ҍ�S�����e���� ��0Sz��g�
�&��'N�5L?�[R%.�)��Y/��5����6m�ڒ���Ĝd��p��,!z5�u&���ی���;�h˅Fn۝�P�?�	U�R���~�i��Lg��x�1��_��iz���y��/��)b�����������V!n)>��x��$;�Թ���꫌��>Y�"KS+���2������U����z�)ǃ�v�6��;	c+Юk���r�k�e}�{�������� ��>�xo����	����2`oE>��"ԩ�ۂWj�$$�%C��L�w��<�:���уe�F�8���DC��D��N���ѷ�'o�:D�.Z;��a�/�G��U(����|��O��!ՠ:Ϸ�����i�D_n���a�/?�~�E�P�~��l�E�әn>�u��8�j�0�2ӛ��1��DB�]��e�!/���\����s��Mug���Җ���c(��A`��qF u�����BT����{��?fG΄*�IX��0F��\�+WB53�ɍ�fuy�&j����X��V�Ƈ?�=J1I�4�궐5Md��bn��
CA�� Q��G��Zb�jԩ��Xj�U�Z�g_2�O	��A�b~��_ޯ����C�"$�ڷ� �H<�/4��EcĦ\�*�9�Ät�˦Y���5Έ�_�Lf9n+Zyߒ��h�!�z���RCW��>޴�'r��U�<���ν'�.�~��5�ު,�0���u6�jb"6�:I���î@k���nj�	,���&OD8�����Y^��r7?��m�2?��5M25˝�E:�3!π�=y�O�m����.sK�E~�`0�����Ib��P��f�۵�x`��Q��K,|��z�c���%W����.Lxd(����ڀ�fT��6�����,0Q4�Eqt��x,�A���a�܏|�~V�d�o��a_|t"x��{���n�߀�Ά&D�#a:r�����N�ц}��rsߤ����:Z�JS�� Yd\�����s!:��K�$e�C�׆6����8͢K��˦�������(A�G{��[zS���	֐�*�{Se7:K>����OG�9=���}�}�8�}�;NX8��~���_r�\��`�^&»0ɮد�h�%�X�l�Ҋ�P�e��nZ��>�qx��=>��~��A@\��ߖo����3��դ!�3e|&�&�YY���vѣ%'	���ǘpܼrSGd�h�)�^�VF�i>���p�V'fXF.2o�f��:���1��Ol�c��Pkl�x7O���t1���B�Y��Vz맞���r!휬�&��B]ju.��p-�X�FF<�$6D"R�Wv��H�GsA�J�N ese�Y��JL+1My��-�B��.�Fi ]��� ��us��օ6|�w@��3`����a�o+�|SDp�=��E�wߍ�p���nv�ȋ0A��Jp!��ST��4q���M!)�r&�2++d5��\sf�V���ԭ#x�s7��?���wf̬��('>��f�^�5?E,ӵR�*,�v���g�R 3<_r��I[d�zK��ן�WYqDb��r3�X)�y=�q�<PS�*���E�8+����9�t���������^���|�U�I�� �d��r	��5�K���F�L���u�F��xs�[.�MH!u6
����p zi�D޺l	�阞�Won`(��/��o}-n����Gw�x˧I��8�D����ފ2fh���kk�@>�K��hLn�C��[#���p��4�������ώ}�M)�z�!|	�R�^��(��J[�����������)�t��.�i���01V����̧���>x�u�S�0#]>C�G�=���8��p�3�Ȯʵ�B���c��D�`�ۊ:�����	b�v��n����s�z��Pg�����d���Mѳ��n�h������şc�X��&�Y��H3�аg�Ek���HDE�l3a7�BGh�'L�A���#d��*��.F�vd�5�sM5F����YK���bo�H��=X�Ѱ�)y�(���.s�N�q���eu5�t�W�\����-l�qj�o��y��ű��������� �XC/Ib�O�R^��Pe<(s8X׷�����^^�\�9���L�R
�B;�?�T�Y�ҍ�k��̶}����E%��Z�F����t Һ��,m��!4u��6��Ñ7��{�7�v=����i\��&	\>D@N��R=�፱1������FQkp����TɦA�^W��ۡk�ⷻ	��p��G��ڧ]���������%�?����|�\E�c$?�t���JLbg�6���-@�>��g714��F��Nc ���6Dʄ���^V�&�)G�� z!���+�d��2�lD��Y�Ͼ�c��z
f̕�J�Ԅ"�`��EU�vZ�T4l�L��Ԯ�tA��9?�j�~�C���%���<Ѿ��|�_�%�N8�V(�vK�M�z�Ѽa��wQ�Q@16mV�:S5`V*�Q����υ���O��nu1��~l�̾��y��!K��Ӯ|1�R
�L�5��J�=[q��/u�����|�d�1�[ ���Ӆf�d�C"��%<��W��|�,:������R��x�����D�U|n�vi�D?���n3��Sa�v[X���NJ� ��x!z:��������6�do�+�5��;�S��U2���ۉ��41�E�
�G��O�s�V�v�!���d���l��
_�`�-�A���5����d�V_�~���αc���	�Y�?g:H�\/�%M�°]7޸V�o{�QȒ�{+�*,��.!���Cx�a"�����#	�G��WՌ[BG�ݧ���]�m<�U�j��Z���j@�3g���|��Fɧ�L4�J(|� ���=_�)����t����������4g3O�4!�اEx�_���� q��Q="<��?���7_XT�p����YR�t��Z��c��D~~}-�ފ�iB�&�O���5N� � B'׈2��1�lKё��M���~O'D��u87��,R�c#��z�s_��3��u ?<�?jo8C�f��$#��T�|�I��m���c�J��v��~w�A�!yDUعSV95�["o?��c��q�_�	�Q�eO'yv������Lv�[��^���]�];ٛdv75�N̦�\�a��Bk�d��
�O�o\����9߾��U~<�53{*y��Z�s-J1|v%���8+��W�ߢ����瓵/����A��[����Eқ�j�9�|�COHM-�/���rֽ�j��r�*4���&�o��vt8C��C�։�k�����"�.��D�)���?���#џ\c������Y��AK�����M椱�'p���o��P������i���G��*��U_�Y�o���>KM�l����͏�k��tgB���_$�.`��ώ�L�x��DP�q�,m�
��H�?{g�-���ۮ�� �G%W�FD��-@D��+�����MQ�l4Sp�{$�v��-��ρ���ќ������@4X������p.I�������I��$�UJ��^H���aozƠ3����]�[��~��f�N�sA��4��s�����@�H
/��^I�����Ak�O	���~
��s�8��2����p�e�4��l��q��d��n�e��~N��${%���E1^��_n���r���F�p��f2���r�G��a$6x�׍C��̠�K�'X!��`
�����g�=��hONѭ =o�t�G:�v՘5�d8�H�ك`���'SK���!Me.7ܛ�"L82��'�6�U���DF�)h��}���N��;{��
�V;��D��IB��W�E�D��`ٔ_L�a��H䤨1�Nx�e�Wߕ�el�|$!���!�O� J�gL��R��n�1�ă[;���n��n_V�;�]6��k�fG��?�y \�U<,\�z����G�G�6lEp5��W�����e����rН���7���8p�|��V�5��X�ꏶ>�i\]Ȗ�6S�4H��)�&� v�;񆢑St�e_P��x�ޘ!I�y�CDO�.U���F������݈������ϭ>�f�loɍ����R�����Ӻ0t��dt�Bu8�ȜI`/�X�ցBJqc��Ji;_�%^v==�1��^h5�T�[8�Eh���g������܌�4������	��es�r���%sJ��@!�@���ӝȕ��0W}��q���Z�s-v=3��[Ћ�-����;�J3G#U.��"����Hc�Z���p샒�n2	g�QT��0[��U�v|���W�B\%�m�4Hj�pV���cۥW4�h�+��� A�Ϟ�n�Q�oߋC���A��Z�zn�Ꮋ��X��N���v�H�0>J�r����B��%P1κM8��穳���9�N�&�bҤ�4��mKO>�ŧ����41���v��/"׌�Ʀ������	R�[���/$��Ȱ2����9�3H��8�p;���Sn�12����;!03�I�͒���Ы��������գ��g^e��:�f5���Jj�Px;M|X�k>7�9�ȴ]��cM���bM|@C�u+��r�l��Ik�km���_Qoh,��q%�O�|e���#�n��p+ӣ�Dg{�rV��HT��J�O����D��ү��=��1���ӷ��s�p��RƋ]��ᕸݻ�}��� 77��3�����&	A��Es�3�Ra���+���F*����.��;�[5s�Xa��oJ�!E@t�+j$o񖇻�+-v��1:��ֵ$fޡ�ھ��OY[�=�F�\Κ�N��h0.�C�l�Fcβ�@+ۏ
�[]Vҫ�{�5�uD�2J���uo/:䰨k�c��9~Lh,�3:��;�0׏q�{���\-��J�f�B����/�ٕ@�o#S|�L���"� �p��-u����r�2��yk�v�ҿ����Y���J��A�8�G��g��zI�t������q���7==_'K��]%Ѐ��0��	1�ź1x�B�'��ۭ�|@�olba𬄒c��|��{�h��H�v�*<2�y�[n>��1�L;�֝D��p}�E��W4ٍ�[`#��}�+�����7,�l(ڊ�q5���7��B�f�
�����V�&TZ2a�k�L�8x��?5��K��ٺ��ŉ`��6���'����+x?y���F������"�⫫+���Kj�p���z�aҞ�~�W�̺þ�k�����7�1�y��I��Y�uK�U8�^�j.�z��U�M�s.d������8݅��ꡋB�5>,�3TG`�7>�$-���PU�K�1�D����rm�3�2%�$��������;��w�?�;�ޢivʑD=���~�IZ�A��$���d�ha�yF4�8�����i�A@ekһp53[��#�~����l�W4Axo���G<���7݅�>F�V"P20���r���$
��y9[qV]�6b�ͧs0�MGLܡq]zq�@8v�$�σ��B��C*�����n �g�*i}�~ ӳZ�װzxu�b�gfb���.8�(��qgb�ޮ�r��Rs|ԑ���^�t��ZRv�����j��E��1��ia�9�_�=u�Ȑqӽ�a��Cq�W*���"��l�OfaS!�5;XO�%G#���M(�ENràG����u��G&Z���1��'5�Y�2��ڧ�D�����6Ew2h2�	ثc�
��S]W�|$Y�1Qb|��U1�{ ���H��9_�8��Q� [̎�c㪂)�+x t����[Ȏ�YR��ج�*����g����,]4S�a�!G\ƛw�(� 
����G���?��Y�£7��7��ާC��������*��V��?I�XFIk���z�dXZ�L�/g���
��̕P�E�amC,)ĕ�@v�S���r
��܀((o塠�w��an]}��6yy@�������Ql�&�؀���io�<�͉��/7�-�g�+	����#��'#��Ir+'��Wi;�4�G�����6��_�٬��zj[�S��ccd��?y�|��ԩVGv���1dCb��kmL��pXG�Xj�|\(��GH�(PK�|@(��JVJn��ޫZ7E���	X�2b�l����)eVn6�S&�hߎ�KY@�!�a׺9%R"XOz�GŬ��c������Q�!�/����� S@鳮#�1������y~���`�=��	sQ��6�� Wa#&F~nʇP��ZP<��ԧԙl)軲W//�j=��L���>X`����㦨���RRv�So�	w��z�7�of��(ѓ$�6���=KT�!{$f���/�9�5�i��u�����Ă�����E��2}1*�Y�A�}��m˷.�V��'<���?� �"�M����~#j�����p�1,�H�"i}N���E�tr�i����[WL���#n�.=N��87�*���R�u��^pO�bw(I�@VV�m�}������g�tQ#pRTK;�:��N3��|'�}��Y0�M*�$ԇ�ꥂ"rǃY�$C���}�ƈ[7橥�IZm���C��ql��A�۲7;:�F^��g�
���ꀲ����n1�O�&)o�'�&���8�G(sA��{���E,�t"N�K�pe�`F�΀�6�6�_j	?R�~~����/��ɴv�9���i���l�q-ۛ9'ț9���"@�#Fy�������#,{�vPk�~��]T�㕯A˖��<`����p����8�b�X!��{	��^�xv
2�Z�l��[]��S G$���0)S;�r�R�IH�o�� ��v�٘l�]���oW��w�w/u���m�ql�c*��P�l8Q����L�?"����������P�8P9M�����ś�L�F�(ɭ7�1�H�����d4E�#Y����V�B^���$��ptt���[?��'!a��ՠ��ަo�%Vhz��hjt�Y$�o�&�g�L	��`�����}��{,RH�أᬀ~ϙ��p �lU`��j�Suv��|MY��Zt2��������޶�b�����R���Zϡ_��z��!#�L�R�}�e ������i&��#�.��y�g��N�"��@{Cw.g�^؉*�(��5�Q�5�.�-c��bHw���U���[�M�ݴW�nؤ��*������nh�T���KW�����2���^�fu�f�'��hy��:�㝧��F.p��s8�xb(B�\-�ٖOy�p~n=��[an:�h�V�C%�� ��w��:"�`X&8b`���$֮ Va��в����[��b��2���� �mǚ����/�HUD䋟#^v
\�n�>G�@�����7pȪ�����v\�����aÏ�A�I��G��]�9��$*�y���A5e��/�"�܊u� ��S�P���f�;��������H5�4�����zcn=�z������v���'Cʥ@̜���V6<8��n�_���G��{�����vz}^
Q]��G7n��pR3�"�KT�5&�,�U�i��:Y��� �0R��~��n��O?B����좄��qU:U�J='�V}�X~op�#��Q-aS��{�Az9+D��{����Af8���+V�� ��Q��#�{9��� 7���K���-D���:M��13z	�����D6�/��	�d-}�<*7#_v�G�!T�H54�y��z|Tt�,���%c����<��x��-�
�*\�n�ݗݗV[��3�-X]Z:V��-W3۪n�.,M=K��Us�AmNi���eC�@���[�W��zm��O:����cu�W� ����RU	�{��CK tɈ���޹���A]��ZFs��7���Q4}~���um���X^0�`;���֡�M4��N_�L	�:��~B[�Uh_�`��&�&�P��ۘ��R���x������>��e׃�"�����Y��"�&����ex��i��])%g"������-�Kٻ����y����|��Ln�U.��u�����V��ya�П��E˧��Fk����2u\7v����5r����aP}�?����թ8i�'P�c*�#JPHh��ْ��]�$A��ן�?�Y�>j�u����~�>"v��5�.)Ѯ=���<�B��HjH����C!�5"Ķ���N��~W�C>�ǉ�6�}�v�7�kΡ�uS>�<��b����ߤp}}=933f�ė ��-��=n�a+�%ra�so��:[顿$^uzi��srU��AVP)�>;�B���Ҿ��H7z9�`��5�{]o1�L��kZ}S��s��+���,�t&�����:�R��V�|����� �a:mw�wv�# i���P(r]�_J �P��1�%���<��g��Ӌ�&O[Yn�B!}C,✩��U��
;y��B�l���)�i�F���Q���$��B�ݧ%�n	k�#�hs��^���΄�,�Ã�1ߩ ��vPp}!����B��X|ײ�[����F��l�������´�v�B+�H����#'�����W�g����8�����1喉�( ����K����U<�]
���j��[����d�QELR� �O��u�f����,��kx�)= ���D0sg�2&_����D"P�,j��]��	DK�n�wS+)_�脟P�pE��FւQ��k��m��0�ιg�$a�`��މħ>��A'�u���*��j���@��Q��nm���*jj��Q��XV�g��x�)��S8�~����,�V���}t������(���/��I��0��<��E��**8$�_(=�?|X^��Y>a��04Fʕ���LF�/L��9���+:{��K�4ZL�*��wAx��8ghH�+�l�k��]E�D�{\:D1�JV�����W:�9F;�]��7�8	c��@U�����'�5�76�H��R�����rG}�ɉ֐<7�s��(R����i̷-�������e�/�OS�����gՃ�M2��R�[��)�1�ǹa��sBe��L,�s�0�ժw!8=a%f/Q�B���y�<�=,/�d׻����L�w|��w,b|K��&=�`]/�Ҷ�)�g�
$�?ٯ�4�u���a_9Gޟ�#�9��ޜݫ��^�-�0��ᱠN��mPN�	hu���;7�.�I,\|��`�%KM7�=Y�"�ͭ��E�1����8�2t���?���i��@e���������״��*������=��(�=�4�N5�.?�.44\�6y�՘�3��Էˇ��/�)��{s�Zq5��v����:��L�"���q�G*I�s�)�&������jbl���PZ=�3�O�v��S�{����DYL�
��<x۝�k��M��!* �7O��i��<b�}�3�B�n?)-8�s ������P�[>��맜�Ay*��s2SC��D�{j+Ѩ������!��d��M�_�+��긇ǳY}�c����~~�׌��x��������i�JUSc�9���6��b-"�q־�=L#'RC������^wZm���x�M
���Nc�F�����ew�"�\��a^-�!=����j�S�APQy��~/��\�"�3�?��{�EK�u5zQ��$b��_���Q$��i����� ��������r1��۪ec!�ޜ�Y?ފy�ΔÚ�jf���#!�?dV؟-���f� ��i�ݛ|��IP��3C~gL�Q^x
�h�9��3��c��_`�LE����J�PL,~�����^Y��E���bq;����w�J��@{��w�� �F�<7S�)`j�
Cd�u�Z���j'0���������y�ͧ�x[w�F���#�
i(�p�ϕ��?�cܧ �@T��;^F��?u���	l1)��s%e������y���ض���ضm۶�6�ض��dc۶�$��W���<�T��s�\��LwO�|z�{�
�[�# 0���KrYe�����	��\��� ���ר���hm������ی�%�i���PV/>��^
��	��ң���ؗ�� ��p*"/!'�U:%1�����pi�Ё@2��ዢfV�n��P��e��Đ�-�;0݇u�XF�vKp�Yi
S�����"�"!y����,%���3_���j+	� ���Nt��7l�z7b��(�ϖ�0��]�iv�ӆ�]�����"*�\���@��BK���Na�|�LΣ�(޴ud37������?LIq^v�Q����%Y�����J�>��DCS�Dp��Sr)^LK� �	���$�'�	?A܈�If����#��	�G�"��T� �7y��C!5۬F+�@Q��k��;���ڵןK�~|c�ty5p�i�ط�^M�\�^�F�z��z"�讔�cᓬD����Ƌ���ǉ���!�����s��A�=A`6�4�|P�t���Sߙ@�����5
����,��)^5�T]h���pz�v ���\g���d2�>~�p���릙�7?,�v�c�ʔ��Hd���#��C�B�Ix��bM�6���O?ռ3.��w����Щ:f��r\Y��e�\�3�[-ǐ\H]��Qk�֜���(]�__�IH<toכ+���Q��T�R��	h�hpSe��YX�;������^h����/S��lV���r%����Nϓ��D����,F^�Od/�"Ƹ3��黬ь,WF	�����H���Vja�bp"��E��z��J��DZ�,�Y��wp���&w��L�#3Q���oZ���q��6�Nr�eJ���1(5n�n�ߤes�̶:�a�����z*��\�p�1ή�}X��D�P�\QjX�1��c���ƶԽ[zHCxgj����4�Ѳ�Z���m�p�Z-�3�[1�n�%"���z���h�f���% f�����֞�0w5]��<H�I$4zPe�w�&��b���H����Z0:�a�/ԈÕ�mD&f�8p;��j�1*[v_oWĜ}G \����.,�]���vA1އd+�x*�h�D�A�Rndwy�̍b��\���wV[�[��ۃ�. 6�������I�E.g�$){I�[�.&}�� ���f)qߥ�>3�(v�VM~�@^R��<"L���y�[�Y}`���Q��]����"i�ʚ�זA�ͯȨlQ˩;*��*��%=���h[n/��$�6u]��S�+��	$}Ɛ��p�H-�H��+;c`1�f1�[铸3!ʭ��i�^+^O&<d��5�:Q��h7y��h��D��~���V�v�ek�w-�G����w�ML:@ȃ����y�\��}IE;��P�����>��vF+��Jp?��r�L#x�X�,V#	�}�t�E���(��6�c_��O��\I�HS�Ꙃp��"ꁉ]x*l�_ڐ#R�fť�jl��d��u�!�>��l�BON�KP��I"6����K��h�"�-rŚ%:�p�~���D���3��y5\WˡNr3� !�E��	oFAq;�x(P�l�;r� ����Xˉur8���'i��A߁�����ȧi2�:9Z�h��ݲ�̺&��<�����_�|'�unp-t�w0^b�7�*8�<
7Jvd�nh�Ky��1~Q5j��~��z�����	�'�5iڒ��G��b�#֚��py=�R(��D�t�RJ&�N�re/��UCd��y�ל�_c�V�o������I]��z�&��;�\�Հ7�`9�#8������J�B�|�Zǵ���Mߖ3C�:��V$�I�
�^�[��ӑ��>�V,�������^�uw���v#���1��I��猡y�ҏ��tKM��MMX�s�X2f��Zdw�¾zw&�Xs�{��x7�=Z�"J`	�a�'f���6�Y����"�؉��͔�ɗ�߇�<z�zȨ�׃�	��h6{���8C,�x���V�;Z||���J]���WN�����+�6��N���쥞�зw��@$BVU��Lǀ��B4��ϖh0�M&r
,\T�t��9�{e�>��3ᆦW@�4�]	?��u���i�=��.��~x��@��ͣ;!O�s�K� �w�ML�`#y��G�uU9�U{bUi��Q3�3J��ڨB7�e/�-@l��N�1/[�Œ��Y
�3��T�>djRO�W*}%{&`_;!�t���X6|��R� q`�a3�nKQP��k5���](�@I�B���f�5K��s@rҨ�B�*����Dv�{xfN����CS@12IWk?M��z��i9�x�T��4������D'`/b��[`k�6�> ����qs���e������%�Xh��#+1
I�ܕ��C:�{���C�v���G�_�]��!P_��^�ig��x�Z����n�k<�(�1�z_�ʟ㧁�3AL pȷ�QJ�<��F][6�����1Q����j�&���:V\#��v�̨Ė�o>��:zw߇1,'W��ǌ�ݍ�u���Ԅ��$�ݚ滑�]��Y`	(��@��FHR^��0!ˬ��)�#Ό����q1b24�4���Q7(�r��H�4�7����&�屘����Z0�#Cj��J�W�m�E�<�ܻ�~�Y���T�о�,~���j�I��!�dS��Xɑ�U�'e(������:����|���������R�\���Ɉ��Q�B,8(T��9�K���$<��%&���K/���� �d�U������ͪ���?~&P��>g�F�(ǲ*��Iv�H�&L�ؠ6|E�œ�x��i���Z�mTcA�!��XBIe�_�S��a?-�y��G�Na��`�1�<�'f�&p�CH�4����� �D'(u6v��a+��_}������z�:�W��"ޛ2��:�Yn��s:�:�o���H-����U7QC*��3 �lYeh܉�L�,D*)��p����b��|d�ܬ���x$D��#	�$����r���b�("N2 J��cۥ���PٓZ�i3[8���F�d6�d ��l��J����%p�a�o��D�R ��Mb�X�%���Ρ�Z�w��PL�z#U��G�}�����i30�����RD��ԣ�� M���o�y%��t�X�o|_V���}E+���������>%+7¾K������o��Q'l�F�ȲD���2`�H�]�F*F��B&�GD����?4�k�6�P�R���v��8�?�B�CBѷz�*��ρ�Q�����%	5�,����
3��W�G�wC���n�]	�|��H��������pw{�M���Z8*Kg/���Y���Kȷ�Jo�K���!��O�� ��2B�?�(��=�"������I�맃��[D��~M�w!�p�7���l�������I<�T���h}�}Q��O��_DfS�÷���J��o}�S0�W;5ͷC]������A����Ai4'﫽���økH��5�V�9U���ؘ�`��e�/Ɠ��Fn$G��mq�{���-��wU���[^�����w���l
E\x� �H����e�>\]�B����4C���.�zz��lE�|;����Wp2�� q��=^*
jAȷ�s���"��ΰi��I��l8u�����Ai���O|��z6|����db�h��M[M��I�U>O�Z��k���e̾�l�����E�#R{��[u1�d�Z��s���Np%�uH�ϳ�Eal��t�5 �$�i;S8a�Rl�>�n)&�ш=�C�- !8�*Y^��}L��|�|�I�Jv��~��w&<[�Y?�H�{�07u�,�6O��gc���}��i!,F����dH���}�Z����E=j�.��y�7}w[ā!�Wf�#++;�AN+�U�?@,BpA�W{M��N�A�߷3���>�Hl> `�
�{���x����r9��~��?}I�|s7�7���kypq7�����]�t}�v������� ̑����,�����Y{�hi|�w�䅏��O�A&ya��tX#� "��E
;����+�@���*���:炙,p3� $��&�+��y��%�h��۝2\�Z|Q���79�FC�����Yd�� ���#�=�y��xg^�I�}O֢�Rc�8�҅�i�U��ϕv//�SA/��kn�.�qww|��[�~F|(�iEg0.o����OZ5;������W�}�*��o?����c�p�� ��ȆY�i��r��$�:�P��{=�Yª1wS�p���Ơ k*��>L�>oF$�c������Lٵ�wm|T�kh15P�cʁ��P@�!��D������;�P��ߖS��H7<X?d,�).n�5�F #���e��9EN^��*�B�[�A�+4✂�+<S�]C��ϰa?)���N����?��Ą!��} !�=sLW�����"��Uֳ�v�y������Ɗ���K5^ն�S�K���?�o>���vIm(?��x1���n����w�]Lt~av��G�۲�-�-��EԷ�z� �,��_�ĸQ\����nVD�n��|Ɔ�̵�3�[���ٗ[�t8����ߵ�6�WS�l\���X�L�;(��U/|&��uku���R9���/}�����k`��Y���}�:?���f�\����u����4������NEt�0'����c����Oo%�N�Ӥ��N�nQ�E���T{�����&e�.t"�^Ox�]���J�e��ߚ4
�.Yci���Р�'�#*j<GP �%��<�Ld�A]�q��)�a�p^��iN�^{�U�����_C#>�FϦ�bH#�T������-"�B�(�O ��  �_���#L34i�L�$s��d��;rQ�P����^\!mT��@�_vNAؘDu�LJ]|���K_E��kd���O����AQ%�@�a��	�ճ1�[��BI�y/���"���mG'�H��Fʧs��B[�c�抳�@ *n�+��s�$�Y��3q�&5�N��%�:��������f��M��w�bYi���b9�$�f�jQN��\�����=�eS����ڛi3��*:vRA���XH�J�Y��4�$)���1��=����1�5sz�}�U�����]a�^��6�~���*3����M�9�g����g����AWco�ܪ�>U��+T� i�-W�ڥ���࢒����Ty;�#�<�[����7E[�<��;�V�䤖���Of&&KL���!x���W����Ċ�/�坉a-��p��ߋn���U��C"6b�{�c���=+���Ņ+0{��M��P�(!K^���M�pك<?7� z
��s�4r�z������
94�5n��Zn�M]w�P�<�A���k�}kX��o	$3�Q�����+DN�+:�"9xz�����4
�j"�Hr�#�����Tw+o�;�c��򺅼�7GS) �:Z��)�ss���ڒȀ9:���"ҙ�9R��T�1�<d)}>�4��sT��v���o9�7�X��S��b�F���SGޙp�G}ȥ@>֖�<��+wxi��Y�Q�&[e����p�S�����.ͱ5�y'��]c�j�9�x7��,3(��
��j���wŪz��v�תc�;��au�2�$x7zH�F>[qK1#LXE����E09�'zyo�l<���HL��^>7Օ��0�1�ݾ/y�8="
��.�=m&.ƒ�[�R�|$���w�/{��_"�2G�~�,b������u���H���'CW�!��OS�j��2S/l~-~���{_X�
q�{S����kL��(����!�j/6=��W�{������C:Y�<@�AH)B?����.�b�	6�G����ػ,�����)��WUOS4EVMŔh��� �	���PN�3�m]	����h��+�S%/Qp�j�H���5	t�P�Q�fvQ)�9��Z�4�3!�A�q�����B�p�j'����2�����&�cCWД�Otuח�y��3������
�1x���@B�i,�
�������Uzs8#���#{ofiN�ɫ<��|&C�˧(!N��p@��:O1����KqT�~�(9ҧ<����,�m���1�5��d��] ����@e��ti�G0j�M>�l�?6�0v�d���O�/+}���
r��0^��'K��^8~���I98��Os�o1�R��m�o��]'M��4`N�O���oI�V�Y瀤�-�A�-b@��SB07�j�%ͤAnD#@��̞�"��&M����"�}RU�PV�3��t�q���'�<W�D?���|���~ۙ��Aߗ������-��%����a���5�E$@�1���*�����-TJG�1�U��+'C/.�E7�ʹ�X8�=�\.R??��rF=1�~̑�P�Z"�g�M���˼zmڱ�kST�w�{苂CI� ����������5�mQ�\�+ȏ,f)	�t����;AŴ���Ibt��D���ٿ�8rr����%�R�t��ڰ��`q�b�ћ�(�<�O6�9i��o��H��M���_}ur �q�h��ÈfA��c��x�����X>��
�,�D�	�V���G�Q�6�Ǉ���`��;L�A�-&h�hd햋_*���m�%��m�*Z.C���QP9�I��C�-��(�.w2��;$���I"�>%���t[T��2���,T�(�%��%8U� �VEk_oS����Z�d�k�CgU~��` I�ߓP�ݽVЃ�/��*ڇzL�����w]��GE�GUU�Q8�q �n^�vF®\�.�η�\��w�9fŧ8��)�0oГ�Z;pu9�z�������8�^A�]?{�M0��6��#gj�.x�SJE"P�3S�Q]�A���j���ܫvS���r�ŧl������`���d�Ω%�F�� ���.�[x�ı��|)���.o)����U���3+CR��h7|!�z�C
�a^��iʰ��IHTFף�aW��a�.3Ɨ��L����W����N5~���$��]���b����~���b�L���0���dӿCXU�ԛ��<�w#|cյ�J^��������A���]N2�S���}3AN����f��K�ަK���:C���H���Wb��Ds�L9���At9�v�=\�Dc!S��zQ�o�y4�qYZ.�A�&V?����&h��F�	}e��0�X��z��JY��8�C�tu}���O$u2��/k	�\L���r\}�C]�X�����f�-��x��M�� �.v�*�n�I'eE
k0ܟ���|'�W3�3x���UB)����>���R��2"Ie�$��0�&C�����5[��x0��:�3�MA;��3�,�X	�+�RՋt֗���6�Ǐ�˷�S%�k�1�~��M��ȷ���磶G��{��/�td�<	��]�p��q��,�X����s��(=�,ڼ��5���7ħ��z��i�ʥ����ߑ5����[^�AT���E{�ւI�Ձ+I��_��Ar�I��
����L��E�ѿ~������.�G(�N�*��S���,𸾐�����6�v�Z���"���{If̷H�$N_��%��|�bX���=�
mU�y�U�
x��ήmA��8����}���~E��������q��A�:i _�O�]���s�j]�1r��zy���^���v5P��T�op5�W�s�?J�bX��{���{5ل�CU�򒅠��Ś'H��|f�����_��{k����3�'��g��b�OB�#���Fd�!�n�������N�K�Q7�q��MR�"����,}9|����SH�F�`7y�Q�!��}%@�E��q�m��v)ܝ�o��[<�eo�"?��Ab7k�3��*Y���X[u��TѠ�x��G\qG�F����G]�ӒpE�|���Rz��TE��w�^���P��{�o��A�fr�|���Al�߾�i��z�g�yz��|�z(����=$3���}k�A*?�7��|���Z�0A �sR	+�����S��$����h�_P��#N�rf"�G2�m�F�+��Ϙ&�5����G~����Q���M����Wl�F�i5��t?I�zv�|�bIJ�i�G��c(Y�.�j�q2ﺆ�M��D�o��g��Ro���>�=$�ͦ޴�^�[�b��Un��'H���m̊+Q��*�vqu$��Q���W�pR��f\��K���X [&B~�T��t�d��d��,e�s�q�&n��>K�;.N��bꠄ��y��J�>˲�	(Y&/7i��jY�}A9�`�Jh="�K��� ;�Z�;�Z����ɋu��ܓ��V7��k���㗏��o��/�#���E�ҋ���Ѩ�ò�
|7�G���S[r���`���D���UM���|ߕ^��Ҏy�����Ej�(!��dh�׀ |�����t
��$D��Ѐ�R/s���71���p��{EH��O���Q��t��K���������R���/s�Z%A�BKI�d�ڹ�q���i�[
-��m� ���(D�nǞR�0pc�����d˝S�5���,��^a�Y��x�P�qAe��=�m(�&ltA_��裫�ے�����V�
��tYju��Xx�
�IX�ź�˒.��Bk��P�MM�r��eU`'m�<(��4Dx|��*k���0W���HcMTb���_vd��DټT���jL��aJ��^y�)�p��������g����Q$�B7g��
�_�wKs��D�I��h4�!��4�m=��n��6m��uq���-��g$d�������̉K�)�ItH�߻7mV�UN���Z��|�"�,<��ff������hv�6�ޑ�ao]W<�	|�Xb��eړ|j���a@h�-���Y��ҿ#.b��<P�4h"���=
=�v��%�$x����si�F����#�{��:�ɬ���x��b����#�?���j>>�~�����r�gO���Q�Fɦ#�y0���vȥǢ&�f���IV�bC�X����2�a�i��q=�W���_ȡ��]�\�1y�[+��T��m��u �[�n�}}��B����h��0U�
5�|��I��?;q���ĵ﵈&�򔜎��UC*y~��I_?%�7~2{��OtAB2�X�Qj �vDC	7�%Rj� .����xޮ�^nWi7�{ҹb�6���C����ke���<���s~1��}̛�e����6u�L�^�'	(�t��Yf�m�[L=����`�L�t['�Z\X]�n�4���5�<ӎ�5�(�`L��w͖?1.��
J7�(�ŵ�ټDH���ۗ@�M��Rs*����E��6��W��0�b(���j�(���5틾��$�iz��%�1�[ȫ��*�-����qO�R��-��Q��<XfQ�,����+��[�Z1�[H�ӌ��=�ޯ��tF׊q����[,3��BM�oJ��v�m��l���Ov�S]�֝eȶh\�	�4yS��Y%y��a����!b��t��5\D�~KI'TW�3T�D��2����#`ڒ�+��v݁�3e�E��.ǰ`y`+�Y���Q��ruw��Ӛn�彿����"B����DM�:03saV��^͖�܅4�W<#�s�$��('��O��v�DU�!�����m��KS0i�"��L��_$C0M5-��sS�w���Ǜ�q�<�[�؀N��QﾏQ��+��wnJ��)��T7��Z4v@iv��,�s�U�+ɔ�2���_��-��By��@H��igVs�����h����Y���z�?j?ڟW��?1�$���v%�pE�Ĝn,�l^w�A��u��G�ƒ�U[bϑ����̀�t��l�>&�2�����?�_V�ڧ���B�T�'F�f9�
I���Q�&A���O��;�
*��e�!��XN��H��y�YP-���oQ�>���f"�CF&�eg�!dNU��OF`��qZ%"؏��G�
͍.:і��kF;UNe�.w'����[� %
.l�_��1A�����ͻ�M�(֧U�hB�ۚ�K�0�+vc�y��-�������7�V����SLef��䌅�{Ad���% �B��u�{7����-���dS1H^��u�Wp�u�q����V���/pB#+z���	�)�*��gF�; &E�_�.׉۴�F@�׾4.*�!�s���+ά*��m�k��R8�[�Ex���ti����̄�$uLA¯#��)0�TݙF)�bID���*eN�)ص�^H6��1J9��(REw�O=fSt=�1�-�Z�rZ�ba�\ixZ.���p�X�cT��(]����D�}'�hS6���`oc�!�E_�c];hT�/��Ha��fq}3a�� |X!�ݸQ[�����q�(y2k�>X��9�X�m?�H9i��w	Q��앷a�R�O���*�����Fʜ���g��7��yAZP���E��bb̓�6�����Ii�ۍ�G���w�OƝU�e>n�	���˲���am�xwr��>���c
{����N�ޯ/	��-E)4U��Aw���6����`h�0=�d|�JL)��_@?}%H	q䇓Cv5����lN�h;(�;���=�L���a�cG���qh5"�'1\���p{U��b�t��
�[Y�b�r>=C*�'g�?�^�j��n�蛵|F��Ct����Dc�����-įU�7����va����I�hr���(n�c�*��K���N���4�z]姙�i����2kn6�u��)�R/�q$wOOpɎw忮0��Xx�nnq�٤�SB�^A���v�X�8��V�V�1��T��h��B�����O����l�j�y�s�*��)�N�7wI�Ri���\�!RR@�N_wz� N�E���{�[1�����������N��U��6�)��M�8D4�2��,č����4n�$C�́�7t,�de�S�W@B}=>e*&�7֜��I0�,�n��O([n��f�Ȋ�]Xv)[��*.�v(���k�'rjϸ��zv����ŵ� ��4R8I�7���`+�&�c���Y?��r``Xe/�^����ǥ�F�sl�d&똧�rce���b���r�jqGiҺ��K@�$�:��W�d��Z��}wuQ,�c���h&,K� 3C��V)��F?�*�n���&��v�R��sG4��=���r��=��=1X��c��,&ߵ��J/���tԨ2_M�*؇Ǚ�	{x����ȝ"}��j�8z��+r�R���`�Q�p���+� %%�\��4VL�)�Η�k$Sh���N���_ˮ��߿��q��a�h��-�(%�@1K%d{����w����Q9af��z�:���g@��щGW����6U�T�:u��<�-�%�\�X���;�}���%2�HyE1���i�O�o��lNG��uKe��&ay�=c8���ª�+���U�l�G����M�`ÎF��_JA7�UuTW9IS^����w���a8{������̭���c��3�P(��W��hx��Ag[+�r�.�K:�������� Dөx�?x��#N��<�l-K��$�="��Q������B)�g�=A��7����$����2�n?�3w/�[د��i��G\P���\���>�\��*��$2!Tl��(��73�3�עL3�I��$��ne���Ryjg���2=s���u�����G�<!�k�����V�\G!nm���� ���N���އE�L��⩪<[ �\�Ɨ��e}�����4�-�DN̤����-U�.�s9"�`P�2&�����z8���IsIՊ�V� ���^�E��K�6�P��A��h]��B8�"��CU����u��i>}��Ƴ�����4�Ѿ��b�����y��x�=vS���F7��;[N)y���E���]�0%�>�=E�v�4�7�o�7�C���p�y3��`S4�HM���G��hlx�xA�6q����zk��d�-P�؈��N��F�Gʜ̤m�9���l�"G��R��TQ�i�vsI&�U��{+�k<��}�i����޳Ηx�p$��v���+��6-
%EJ�9�5��]�g�о@,���x�3���������Q��j^(��� ��B̸�fp寵��*lIFL"�S��r��3
��
veh��{_+�K�F��帞h#��1;���{���ƙ�*z��5�%;8T����N�^ �(J��i*Ӏ�<�.9�Ȱ뉝r@ ��2PE'�q������bE�I�������)F�W��	2��t����i��V�� q2�|ը�|�����c����ԟ�Nt��h�x�����N:���7���q]*޿{��i>UL�NT5g��ҁ���Oك���u)=0_+MuQAI��9��V��?6D;�ӧ�DL(K\%��_ӛ����ո���X�	�B���ʾ����J��oS�d&/[/�0@"b�ӕDpz-5\�f�f��E�/.vG�H��mP�9�����O<q�iuݲ�)z��̣�V|z�A���q�kݴ�?�р�=���m�j���bz7܏S#>ѽ���n�$u����F�N�f���4jh:��ܯ������Q��3f�ܐ������m2Z���!�A�j$D�pzڈ*���ԅ���`�!�ӹ�j��jPsE�?Q������)lD���X��k~�@���b���飵P�Ѝ��Ș����*�RM|b%;�	h,��[}���ُ~6n�]N�n���m(�![5�E룡�bVc���oRGK���"�ŋ
l�ՏN���ߦV^�z��o�Y�?��V8g�&s��ސʑ��Ҡ���[����Σ�b��+/����2��ϜaȾ�F��Þ?Ѐs'ќ���,�]�d�%��R5�ț>g�	0��a�](R�c�J&��=�oH�h���qzW��$�J�=�L?������2�#�Q�K}��V�n�e��}}Dk�� ��e5rq ��e�z�n���^��D�*!���	(����,���2G��ӧ˸\�:���jዳu,�.���(Q}����ˀ�Oس*ICбn�6��}����/^9�!V��|=n�C��Y�CGf�G�"��ux)��!P^c�	{�l�~��RJ�X �k_NO��p����3L*���E��K���:0���CX�h����L1D���b��)m��`o7L4E4�y@��d�F9���V������Ў������8���rmV
��hp8'��Ҷ��j����5u�v~Vܟ<v9��VC11���g�F����9YmrOFM�9�󵩫σA=�"H!v���fF��CE�#�x<�|��g,�P812��l�4=ʚ��&�o��W��e�ǫ'��-�P��K�-�����?��5d�޼�pgt(�#э�Ő��	�4��6�a���1�rCMHG"�����]���V_� �_�����z>`�<���-����E��e�TNgP����%��	�%�O�n��ԉ�G*��k�{YK�
�;��6�dZ�pC�n{*z)B�C*^�eU%��p4~�k�)*�mj}{���~�k�1V6,�+�YL"@x�|�C$ SXӉ.�<�P2�_ b����Z]�s���ٞQc��������r�N�� �]��X������ey���A��=����փ�Ǹ��ceO��)� ax�o��'|�]�戤�j����`�G���I�u�&�=8J���F���!f2�%y�?ܥO8Ov���xu��"Hy�M�b�<?�ע���ɤ$�^�BՄ�	iG�ƛ�6���O|�!@�jW]�+����]$�_�_���$�%_7�PǑp�UH"(<s�^��<���-�6��)�e���	o�A$u�3��-�\��p$xv�-��C�4�~��x{ĕh&���u��D� �*5%�y��8��ȣ��e��M�4Q�݊l_�����w�˚8$�64?ب���k�t�Ѻ��Zr�s��b��ꨏ@��\�}�~����\�[��3��a���$���v���Lǚ�7@a5U��[�[�Dr�J���i�ߞ3���yY5 1�`^G��y�|py.F� �^��[�4/=sOV�f[]-~vI�ƞK�B^�П.k�(��[D_�!sc�i��ݜQ��
������|��_j�C��w+�@�γ+�i�>����E@��z�BD��f��w���.�=��4�ܐ���w���gN�*0���j���D�A|̹g܀(G��{?�JŶI�2���j~,[��]/^��5~�~qh�N�J�}���	Ȉ�,��&n�H${�/��JX�Uj�@���5�w�2+RSV�s���$.PҢ;]�'�mDR(V��_R���us�|�}er�uz��b6��.�%��#êipU�!D��w�z`��f��i���{��@#bs3���I?������+�F�*�p)5/*��.o�<��U��X��d<�� �i��7��ȏ)yr��N�9�6���#!I���n�S���;_��J�'��gz��&��?��Q?�[�����l�H�5t�N&§����r���e�Ӂ�3�}.n_W.�y��!�N9N�
�<�o�ϖaS�ק�3G"����F�����k�jL�������0P��mr)� <�,��x���9E�
��Hp�Œ�U3x�2s��������$������	�o��j��2MqL19"F�%k���C皢�5�v�9�m�Q�%[!��4A�r*{��@�`j����>N�~��S�ޙBƀ?����6��0"�_p�������5�y�L�U��2ߌ�^?{��5�Mbg��Өվ��{���u@���]���ֵm�<_O	M_�}�Y����irM@�(��Ѣ��oa���/�;��C8�R߿!�o�;���K�h�5�Ԥb���7������1ڸC+��H/��~NTi����~�l{�khg��K��^d��	��ˋX<�g����G�����.�[��l����
���9A�����2�O�V�����-P��쬙j{����~&T�Z�A���9�K�[JT�^)@eG�`� ����w3�w��Ĝ?�k0Ҏ���:%A�ݟ��	Z�"������^�!u�v45?<*Tq������ʺ�}ɉ7��ZD"�y��X�t�'O���.�4p���2�(�'��6�9��	8��E૭
u�U��@����PT��d\��dqG�ͽh؄M��+�@h~�Pq�F��ph8�R,W�k3�,!xrH�|ڂ"<�瑑� �� ������ t^{�C'/;ڸ���������=u�@�f�N���k$|,j-���P6�ym���>��
�h���:����7a�S��*�u{ⱆ����{u_���� 9�>S7�)k��0vJ��1n*���>6�/�ք�Hs�t`��5�XPY�k�V�S	�[����w��W���i.��PX�A��G�->8�p�%Я�����)i��q�Y� B��׋[��l��x�pGVg��//����;�+#�(��a];��S[�����8�nA�iHr�B��t?,s�A&�d��O�E�����e����p)�R���ƇHp�<{���)p<�2��ݮ�Od��(�V��݂���^�.^O����U�i�H��G��O���U<�v����Z�'�Hص��TUE���h��.�����4tgϓU��}�!��X�ƛMȢ���&�"������S��kC8ȗ<��;$���>����d���2h��tM;N,��e�ё�B��#�����ՁA�##���Z/�+��<�y���N���6���wQ�y�O���-�>�kt���>�:��`A@�����@I����И^�/K���.��k͗��$��.&ܱCӅ �ϧm��Gk�9EU�Xw��.׭fG��~�sX���`t6[�w�ZQxrA9����ޥy�or��_�����(���Ȩ�J�!"g���������;�e!%�{�	�r��Z�����k�@[1QO�/�%-���M��X곞]TK��RS���ؓ7A������:Ɖ[�ec[Tg��r2��.��R�B��qb���`�C�f6��nm�!]�}�@��Ҫ6f�gS�u\����EP�����j���;�FY�ã�C��D$66��3J������t,�x�'�����co���s'�7�����ai��'W+F]����-�oJ=>��[��^Sa�v���?����`�G���e�����:��h.k�5�n�dMKR�HV�(
p;|ȑm��T���AV��"���C��6��3-R�".�H} `L�PP�f0�
��"��R<�
[����O��f�2�8�/����.[�,VQa%�@�����Eph��KX�O�޴�������a�3i�el۶m;�ضm۶͍m�����ضO��qr�w��QUOW5.<A�v��@@w���W���_:7&�1�"�VjRdhʗ4s����ט�T�j��O��u����K8Ë�P��^�x�u�FH+���lY�� �8ד�MMf��x��w�:nU��Jm��@z�2��0Lc��g�� غuw
�}�3����J$7����區�YqE���p`�T�	�ۢM�KNC;0��Ậ���</_K��'�y}h2��@��l�] xhDA6���*��CJ��wHDH���`Ԫ��VԢ�>�"��5�N�]7.�W�vtk*�����̪*��م����b�����_����k�N���n<=��|�m�jC&J��W��yܴ	��e.t�b�\X]Я5�*U��U��xdp���jm��S+��m h.�Tf��
�k�A��IX!�LCM�e��	����
��Pq �9���>Wqώޅ�H��"X����!#���`�<W�ё����&CHڅG���6�d1#�7U�B�#����-Al����kq�݃��{	�큩,�����![M���~����F?����*4���ti�@"v�z}r���Q��~H0T���>��ajɢ���t۫dSR��ԡ�@���wO�~N��w�Y��E��?���F<�71	 в���=�a�SR"��,I<���봶��'��"�B���dK��9�Ý˪�h�j����E�@&�e�*��x�43>@!tŎ��a�Gb��Z. �^�~J2Ӻ{GJ��,��Zy]z���������\�xT[@����k��*��.�ip�@ �4/��|Qk��zw[9��+��u��Q8z6<h�U���f�dP3x� E
2�
,��cL��{Ug�,�RB��+����1��>��?I�3T��=�u�zJ9ϵg����=��i
���6�4K�ï"��a�L�4^����'Z�*�"�{o�?�=}hX
�����Ԩ�#���$�|%#��]k/�����kt�Gnw��1�˥S�55Zb(h�2���q1��r��N�����H��>�0����"\!���	Q�Gm�1$8fv�e����������#kw�_��]��\����j��n
��x�dz�i����.�w��(Z�S����y�&�A��/��@�Z ��'����q�9�!_�&)�"��M7V�e#-1Vԟ����@����0�^�Z�!�|o�Zu�;���j
-
:� )3uC�Pe�NN����	~U6�7p���׃�+�Z�����-Mȑڤ�1�����g3��Ϥđ��t�?;��@_46)v������:u�~�\	TT ��xDP�ˀb����)*h �)�J���>>������:��\�@�����V��U̘��Sx3[ɖG>�ɦ>㤠�/��#�bӘ�l��ZID�û�1==:�@n�]Puv����ڥ�A�N�ֶM��ܖ�h`;���`we?���2��H�����dؐ����~���W��yx�m�9{2����kFe☛�V-Uǔ�Hzg�knk����:�VtB|5���{���.�F�ʾ�I�5m@ 65�YI�Ή�D��y��@ ��|E 2E[m-�)��0F��˴��v@����X�%��R�)Pޔ�����L����-�H|rJ"�;N&���nY�e�,�N��7��������S7ޥA}�>W�%P�`�t����8g֖n~�Y�Um̂'NJ�}#�J.iW� 'rv�ς[Id{^Bl"dȴT�He~�.& B1P��e0=.�jo������
�s�<j������e�&��Q�t�u��1/_�w�Q������GId����K�c�����܀���b��)����!'F��޶�?���$;��V���Jmo�g6�j�qҟJ�BI�8�<I)��ǡ�u>�S�Z�~�H~>A};0��aNMf��u�黟Mc;O�����#;�L\n.G:R_�Ň_*�J,����fҨ&;���q�a��`mnh���6'&�����oA�Y�-P)�.¨m6e����ܾ�t�hP�0���î<�^���u��1�ޖܽ��xWl�NXeD�g���J�h�qsi�郏����L�Mc^!�m����X�_$l�)�յKs�EVe5�����ix���7�=�/y��kY����>YN��]�Gﯦӯ��O�k���Ӿ�7�D�^\"1�� ��_�A`Q�T9��L]+>��\�����T��E��WvSf��H����R��ZjW��?�[x�34�Gy�4V�w�|{*�q"�� ]h@T@����)���y���PAe|^)��<.�+B�C��ߛ��
|�_�5���x��Z�bU����N����9�*q��R�]85��D�in쇵����+a���#s��A�R�f�Z��0�����,�|�a�h!=�~g�%"�C�����נ��]��Pf~U�J���o	T�s&K5upVg���Fw���_�l�]�#8b ��R��'�^��K�7��^a�wd?�-xr�c�4,�Z�7�B��#��˓�6]5�M�����{@{��,)������EY��]��n���t%�O]2��R�alb�)����j�1���I�Y��l&���*ܒBh��lQ�ru��Mw_��:_�q~�2���|�g]Իfngڒ,��^�ۣv�N�,�gBu��+���i�9Sw>Y|���5�!ojȆU��ऊ&�pP�<���߰{���:e�RǜCB�<Hm#X1b�R�����S�`����G8�i7`z�
���NhN(�#����L�I=�/���Ǒ���=�w�Z����'�x^N?��'{5��w^�?*7S���Fc����u�{��Z��iM�/aL�(Oȉ�#j��)xyє:c�ub#4���E,F���?n
ʺP�|2��1t�a��cy��
 ����`��TA���BU%���Y�ͮ���Qg���G�$9H
Qi�`�y�"X��j���%�jU][�_x��R�M>ݴ������m��(֞ɔ�:gC��5���j�`�nK�b�s����iI�Xo��D���̂TǬ���~�MX�L���Y���B>]T�f���!���՚5��F�����(k.�����}�v���V�?L*k����k�9RYC�W�Ky �o^�"]��O\�
Y�e'���tŭ�zb��h��x̑6؆��C��`$L��@�N7`�f&C���p��E���0�s�`5�q�"�@�Sn:���#t��j6ӶćL���Ó&VJ��S#U�<��p����*(��y7�~��r�L`N��Es��o{+`�4\�tw��Y��G-��vDRd���k����i���5��/�t����&أ:|ӥ�r�y'�{����ПY'��?:�L�� n��0�A%������<�o_C��Dp"`�;��'��l 	��/����	u��^u=�8�J=Z;?{��4{rJ!���h8�4�5OΘy1r&���ւ��|{W[�q7tTx��Z'� m9��߯>��th�l^���	GT~/��� @��YYQG�u���o�m{�J{C�B�Qi���1}���䌃�|�+��R[�=|��'�TI���55�8zR��D>�񎒳j(t���k�Y�'�Tt�s�Hs���������F����&1֒�����8!��m��!;�/�iY"�?%�^F�	��O���IcZ&<5�������MG��A��k��ࣖ*�o��g8�拄n(o:*����7A� ���$�n.~��޲S��g�+�ȃ�mk�!F1�s#���m~m�w��pvE���S<�NJ8���,���2�5G)$,�pW�usB�(NH2��u������yM��Au*�h��U���j�	3A��O�S-��u������d����4� ��Ӝ��K����r
��Џ��(�S� o�*��g �۸P���u1/��?ONV��DϤ�u�E6�[��3��B��fC����Б����'�����!I+���if�13h[霅�b�1�O�(�N[:k����J��ĀF�
�[����0��E��D?��D��cv�k!b�H����`C���E�BD���F}E��8班�:��~�*j��*l�i���M����Ci�	 �4Ј%��AV0V�?��cܞ5&Sԗ^���%���z�Ƨ�F�A����3�$�B��L�� 䖁ǻ� V��O ���Y��8��x�)wmz���<�Ln4|��m���Aq��0.������C�g��Z���$
�,�	��}����O��--�*��D��8����%.��+i�u4���|V�;��f��iɆ�R
�HپS���\C�x�$�#7�-���?�:	Z*?�T�1��zxCڰU������&�x����z�,H�|��#`��k߱r.��4����+�qI�����8�CGʅL���l��&d�T����am\������0������2=�ʳC��WM
MҜ����v��;s��l@���w��p��J����*���2-gQP�HK�>��Ү*�M�S)��xr�hf��&� ��ݣ.:�8*?z�4L��@O�u$%O�fR*��nڌ�}%1��d-'i<2Ĥc���u��
�x�������N�!�6�F��n���ނ���M7)����żu&�K�^�nq)@��V��1����ʉ�<\q�E�!��C���vi��q����Z�DF�9���uS&W	$@d]=��������S�|,]V�gCf�Ƿv��?�>.��.�E-o��0��y�P��!�Z�c��T��Ѧ�2��	 $���ȧu���$)�d�2���մɠ"�UR�%��?�YN�s0|�y�v���RT����˪��M`�Y|,�G"g�뤐q[S8����i֦[��&�(
��7��_��&�ח6C,4y�.�h�����m3.�G߮q̩g�r-Hx�S�����Z&���n��(�Bf�*�-@�	f赵/�k��/���R�']�@�ѩ������{ھl>]��k�4���=!?��|0u̬��Oo����-��m;e�MF����z��	��ߜP�o��H�U�r���ȡAM%<�
"�]�q�_ki�H���$%q���
q�]1�|Y}��>���Fp��0�v��-�aO���No#`!���a�k�~����k~,�H1���9���)�z���Z��e!����/�$��uuweP
�����6���3�����3$ ����5E3R�L%��t	��FN��ɠ�ٸ�"������M��!��'���r�3M�� Nb�Y¤ض�?����0�Q�(���K�p-#ASzϋ5\��ߨ<�|I���j�J=�=����H����[��r�v<^���m�z����9B�9,��R�٘>J�A�f���jT�GSү ���`H���:%l|px�p�ԩ�(�-n�F��3}\�-� �9����Gr�J���a!�2?}VЊ=Ԁ��6&¢m)��0�%Q�<T��.=ֹw!V[Y��0����Ħ��I݀:v���ãaK� w���	d.�bz8'IQ���G?lU-�� &��{ا�\U�k�d��5nC��(��q�g��0�e��2��[L�{.������/��;I�{� �x'�benK�1'e�#�S{T���_�Y����ڝ���6KB�|LA���#)��I=���N�Rn��`�����'�,Ψ�cIq��V������{���8��@� �b�Ĉ���ϙ�粳��.5������	�)S�Þ��ٚ2 P<ya* g��P�N��P�'@w�9����~�,���!��5���Q�Lp*��d��R�	���h�?��l��*_cg�)jeY��5˸�ui^���%�LUd�D '�Lź���3�h C�|�P?�:��E��6����BIp3ư�䳻L2X�8�SM2IM�R<$Q�6��E8��#������(��;k��n=:���k+��nD����Un&�VMDrݘ؁�]������k��p�"w��n�����oO�6d������_՟���siG��D<g�k�өN���1_l�(0�|���!�S��&�����'¨�h[�PeK��*	/�D�u����3hD[|�B	y��B������b��)����N_1��[w��R���(���`Ч�l����V��S*4|��t��g�+�B���,�2G>�7[p�KK��-�b��v��ڃN���50��!���ȵ|��e$�`��ć{
�Oo>��_-���;m�5��Ez5�@"9���2���!�2d�!��fs�%�{���ۋk����l�b�;�jn"� ��?��O��fw��4?�|I�fD���HY& D��6aX�f�*U� ���ٳ
��k�rT.����S�/��8+���=X��}�t�*r�X-����TV��eO�r[�<ˏOO���緑Q��5	�iE.��\�یpgT��Ӌ:j1���G�K+����NT^Y��܏�g�n��Q��w��E&a�_�d�F�(��GӨ6�u���>}_d�-�o�@�6�J��D{P��8����� �
�W��'����>�V`�O��<q����#j	d�!���\�{@u������e�l��z�����6��	>iL��e��Y= *�s�������N�m�钀`������j�/v���$��FQB��fN�`n��e�duygJ�{(;����h�fޏt{��2.����_$���jΠ|��x�����Hf(�kǼe<�S��9��s��a��Fd�VΑ�� iӡ�ح�*HR��"�|�Л��y���`qꜹ{�H��ZCm���߂�?�v���a�������ry�#ď��%�W�9���9���~�m{�#t] HftE�4o,ԯ����o�~<o�|���~��3_��r���(Fw�I�2��q��	 ���d�B�3�f���y���y�NR���fse�]򋲺��q���;�_W����H?�h"�05h!���������Ǽ�
}�����˺�Aj�q�Xc�>ׅfhqu)�f����R��_�\�2�x��b?y���,Ӵ�u�!Ad$�4�����]lP��*h�0|�>��t+w���l�>^uf�R��=��J��A4dL���T���R��5�����vh�³�+ī*�m2e�V�$]�Ic	�q�a6W�cA�^I���n^�yM�!�� z��r�< �_��<���1~c��%l��!�"�W�?������(Nq��g�v2z�]|2���ʀ�G^XNv���w�����~��h����=H��{�-� �W(�x�^�ۗ�b4J,�w�H&6�-��Քғf7��J�@ ��4�#H⛭�>%%`������x���`J|n��+�+B���^��۞sO�W���$�ݬ�'1ށ((���NY=N�ɰc~��
e���#�{yDL�9�,iq���E~����}��`��l�&����4:�0�R�(DK��g~#:e�����p�ԫ8��E��?����4$������g���#DzMX�a���`���_��d� j�� ����lY?�C���>~]��-��t�k�<]#�:���E��7B_���B܅;��l�'�~��9��C����2W��t��N��@�}�-�"���Ϝ
�O�P �6�@5I��q� �=�α�OE���ս|TZ���(��s�>[�9*L������tE�B�#��B��� ���H�%fO#\�%��֦ک�a@�1� �I��A4���aF5���c&�L<�>���{��?]�N$gB�6� X)����]�B�5z,���t�v^�*GÀ�LRD�6�Q����;��Y�"�X $���#�c�� �+�?J�T"�|�_��_ܘ�f�>}���-�-͢��ҍ�����Hnϖ�$d���O�E��O�i�Wj�MǥV9y~��FZ(N'�'����S%d�pN�<E�R|��y���љ�f�S�_r�[�%�*��*TC4�&���
œ��
���v�5ɭ|ۅ���Z�td(Wirp����q4_
�A��c�ǘ�%a��ƶr�>Utl�|
�_���i+�?�9��&�g���D��%~���W�j>�Btφ�s�S����&�2���s���D����r;�4b�͉A�.K�x��Y��+,N��v��ϵ����E�k�#�$~B"��������'Q���n��2:�_�V�s�A��P�`��2E���M_T+�1K�����9yep�:�J���4k'�\��,�E���Y��eX�����:*�>H*Je�'7k[��X_�K�vR[��۶C���L	O���ɷ)�f���Qz��ѕ&�ʄ�Y�ҫX�� �A��=��4����'��6��Q�d��S�O���LQ�8<�z¯}��P�=`��lF�ˣ[+��U�o�!�"��^��������T3���C�����^�nEj����J&y�L���v`Ѫ�%�X�P}i�$�Df���pq�;y��ٕ�F�xJZ�;w�b8I{���Ł��d�>�_p�"A�U�Cҟ�8%���V��<9LK&8��JWή�H�n�S���H(�����"q>�q�L��a��@]�Ƭ�#���-��5ax��	�9�W�7�X��p&?��_��e�\1@o�����{�#j��.~�t�K�{�Kl'���7��`-nm{�9��_�%�n�ߨn�������ٌ(5��1��&��p!���R-uW'����M����o;��j;fF���"��Lp	K)hT��@�a/��(� �puS����1���j�Y���N�O߈f����'����vfaa�+9~���Mf@�x� �/ FXNH���``�}�ClD��x�'�{��T�8�GGe^���T`b��q��+}�����m��Q��B�U��xM�Zc�u�\Tkl���Rhd����o���R��ɦ{e.|�����B��׬P��7+�~U�@W�͑�O:��C�
~�q"�K5~̓ΐ�l��0z_�_&��/.�Q�!~tiU�-;��_ �F��ĳ�z�t�}��"��y_�f	E�˔�i�w�K��ݢ*<��8x�ٞ�i�_yP�/�Ȩ�L���gd��!��X�Xg��&g	�a����|�� ��QȌyb���/�AR��ǻ��T{�# ���@k�x�w�*����&��������}���y1�T�/p��⬣l��H�#Ҧ઀Y.�cD��������W�V�A�x�%l��RE:��~L�Ya�}��U�=s���9|$����� 5�&g��H󲂂o��/�b�a�ϕ%���}��H�����- ��~'����*LF��������6f�����h�h~>s�I�sϓnX����,�#'[cVΪ��}�����+A�:}o'��N	t���z��nik�Te{��g��x���Yk(�Ɗ�)�Q�M�Q/w�tp���k/�J5�%a/�/n�'��d=\>j���Y��띠b%X��T���p��I)JljA<֎��Y�8���l�e7�l��qGH�H"�|���-5�7�!fe5	�5��/ءi�����A�t����o�;�7q����͟�����S�j|^Th������L ��\���-��K�x�9�OUq[���oq[Z�	�"���ߩklЦ�_:�����C��R����9�Ju}O��;�JMl�%������pVvk���Th/�U��f�UG���
�&�n�� �,��@M�:J����"k*��e�,�E`o�X����S��:��'����eT�����m˼���u��mݷ�Ղ�G}8#]���1h{���C�>~!�B[��x�E"m�%>[llt�]=��S��@p�W��ϗb̐B����G�F���1l!�S�A�aX`�H"��M2��?m=J��º}�����/n���='/�r0�V$�#oq(0��r,$i��LGlE#������.q���=����F>��,6�0f?�ѮF2�Gĺs�&�?3߱�&��D\Mـ�1��V�.R���T�C�,�B�H�ڇS����u��R	=7�*��$2'�W�X�9���D	`�hD���M���������5U��"A���:dL<���Z�z]/���JMI���
k[���9����� $ݝ� �|p�"dQ���P4[{o�7U�Tx�f�N ~A���)�L�{ݖy^�y�BW�K��Ft����=�� ��FXGlk?�b�Z��K�A���Y?n����������Y�;�c�go!�$�)���Jja�wD���X�������+����b��&1�����t�U���.~�bR3��ʔ7�\3<ɢ���ɞ-�r��kT�y��Ǭ�w��az��d�"����]yy�7v����b��۽��K`�Dz��f�Bc}��v�*���.�p'_XL@!�&a�k���"ؓ���FR�7E��t��G��ѶѶ`!ߟc����n>AY[G�LMG�%�`����j�2�u��G�[�N����� ��E�y��"hd"��WV�ES�f�肩h|=⡅,=��d]M��>W�l��e����X����қ��)�"��C$��	&X��b�t�D}�oB.��z���L��݀6���UBF:��^ay/��|$B�咃��K!�[�l��:�Z�W�dQaRB|vXۀ4L�tV��T��	��P1"��IYeGx扡d�����Vl-y����X8��C;@W8ҘrƩA����+�NbjJ���#8��[֌�^l昡v�;�O�)T��3���x������@_j�=��uv�7�J�Yi.�	���PC����Gg�ln�H<X�yoSР=3cb�%��lY�N��2�A!��>J�����#4ܚ1��T�RH|����lra%���O�7������m�TN���ח� ]:�j�$$�~?IF!�%ò�KZkw,��V	H�f�7#�6z���<�|3�����	y�	���bP�DQ�ۮ{�L�AW��l�Q\�b������n�5I������{��� �5��X.Ŗ�i�}>�蹛�]VU��mf�8���ה�q�"����07Ŋf~�6O��+q�;{�{z&��">�)�=Qv��ȓك�C$�??��4�R�MHO�c�`��&"Fj�ЧE�^����B آL�8.¢�g�,��^3oCO��軒L� N�| ��`ы�nʙU��K�脭�g.����P�J ƖW�)|Z��Aԋ�r��<�4萣�-	%�~�_C����~��ȧp����m���鷗ws)���ZRy�ߞ�����U�3,��tYݷe��a��/M���*��eT�f`x��H�y��/�f�uè���*�َ�4���2̈́�q��z�E�\w�gd�s�2�lԭ-�Z)ܱk���5pU���f���t����5�~ǣ;R"a`C*��qb��v��W���p�*���k1�Vo.���1�5�U��9�DTfo��9���A�kU���kmhQ%[����ӾR㑱?{lj�j`5�u���e<ݑk�|��/bk�_e�ɋ�7a!�}�K�9���	!բ$C��kz������
E�x�����\���?���Rׂ�3l��
z�S����d�wК��T]l��߱��(ÆC/Emu��O��^q�2�0{�
�FM��:�܂rv�j��=8 ���G͠�;�I�Z�Z���

��_Cj�{�w/�?s:��w��k�J���p��VO�Pl�TL��+k^��c������\���F|�ê3^�]n�'�_J�⢇�i'�	�[;�?(^�.vܹ��0<̠�į�
�)>у;h��~��t�}�6���ףġw�6NG�  Z���lQ~���V�.!��fr|<؞	�CW��s8��8�~
FB/�]?,�g�pa�r��0����Vt���
/�}a�;�W��U-K����;8��w���?�#��:�qP͇��dZO�)��nM^�^ك��nllA%\���t�P/���;�֕�oZD?.
?�H�2��Y��Ȩ^HKg5/��.����H����`�׽ɞ=�y�,R���l��ag֕�b}�pN��j���d�n*�'���iS�����W缹�޷��:y�?�c(H4�I����ge��E؏���r��K~�#�IקةD̦G|O�����˛\�x��^�Z�n����&F6�$%1�evj�¦[���Cq5�Q��p������x�\�z^�����",m�d�P=9�+��V�4"�+5/u4��&��O15? �$�� ����G�����c/�G����DW��� #�%�Җ����ӢѼ��ް�jb��X���6aOc& ���K��~&dd�����v��4�b[�+l��qX�X��0�g� �nm6i����J�e~v��00��ز�E��������P<�a5�0u�r����K8r�x���H#�����s�,�JJ>�	�|/�U�ʚ��*Fոo\v`����s��z&�R�#L�����+|w�S �Ƴrâ؇�S�e)i#�s���q��u�.�ϻb�o�1����_�y���@%b�ҞA�3� �b`R���;J��A  ��8xz/Q��W[��j��h��S����Ui!�6��ruv Ը��
�/�����uV��������UB�*A��`ԭ�/i��z�㫕:_�(�4(�$�"U2�
u����VkЪ�*���<�7�⦋+]�Jr��X���bt	��X�-
�K�����ɉ%�H����T���cG�5\U�潊���'\ -�1�ϯ*׬�s1���ڋ[_�s�3,�h�=S,a�
ĳK����1����F�uMFg�O�?; �8���	� �p$&��R7h���Fd�~Qn܉��讶�\4g8���zU	j�G�Ea��NK֚x����i��#}
[��[P����G�x	�kB����u�s��}(��T�o��t~G��S�Y��֬��z�;���Y�!b"4�+c�5]�_�xm�ݙ�~��I��9y�pN�� �.��y�>�qZ�c\���!��6�Zh()�hD���u����G��u�8�c��_��x�:i7�/��6^�e��B�a㐀�{��Kc���"�<�=��s��;jw��{�Y[��
,]�h�n����:����ןo����EAz�Z��@�`w���;GjX�L+�� �B�x����?ns�{k40#�{���oۿ�Zё��q�D,y���-����>~���nh��Ŗ�RӖO~�u%M���8F.��P?X�D���n�E�ye]��e���c�"�ޓP�
:�4�,�=6��\L�/�nׄ�����cS�֮:$��]"�\^�܄I�|e��ϊ3��ܦ2�*��Y!��:J���s1o����������c#�"Z{]���4o�=�|�zZS��La1�N��*�bS�̒�x�t��<��,�^'�����(ų�k�t�I;�(�8U��oE��>-[h��J����a�!+���3>0%3��o�}��M*Wc1��L�5��>b0��YO7J�A4Q*�l���,ō���m�:<�vMh��iCA&������a-! ��x����k ��l���Ɍ�*7��p���Wg7�2N��Ɨ�����V����PT,�)P�� UJ_���1U��|O��p��=z�qD ��H!z�m��i1�HyE��?����3�E��l�x�g�鯌�6o�❢�����@ƞ�Y#�
R��]��Q�&lI�������8�N����9�w�%T�4E&U�0P��Sn��\�C���O�
l�6ޓ���35�Î���������4����1$��!�W��a�>�T��y�u��>���e-;��"���S #���p��Ɇ�O-��S��#��彛=c���Ͽ״����0�I��VE��T���`,���-�e�:ybg-��/�XWn�]�,���nD@DL�"�1����榾 ��c*zO�j���R�!-� ��:������=��sqi��`�n�4����	����`�;�Y�w��"6���
5��y���V��Qw0����H���q9=�SS���G@�O�#���@6��˸�_��[���\6�9���D_�u�=!�P	�ܰ/ns$���s��w��!�2�h���9�Ɵ|@�M�'6���R���E͓��ͽ��Z�.|�����'�MĨGx���R��I������Uj��I���O��l۵�r��q%s�d(�>O�r����0��|���i6k%F��c��*鲙�X�!��Pz2���XE�9�~���Ŀ���k�,��t��l�qe��k���ގT#������4���v����^��+�$���ګ�\��+Y��('VE��jj�Ҵ���rqv�.r��<d%&��9��	��\�ltr�7�������^���vp�`�F�1QP���s�y����b�#�c��2G;¥-�56��φ����d�&�DF2�yx�| �P��ռy�D��{�����[�E��	�9���q����g��N�i�T|�-�3lx�oS�v"����^[�����j������I�S���;o�M����|�\�����J-�2�k��7�>�������O���!OC��3���C�M�^�95FG���Un��[\�W@����H�(��3�J�?��:��+�'>�ck�R����R^�>r ���#;w����*�f@@�Y*�iQ,��t�Pd��`�c'	ԻU&$������u��]��	X�k�kK��E��lħo	;S�K~�	��X���n�`��ʋ�Ƿ���ėk$��w[�ő�DGˊ���T�ỳ=�X�&�} y �t:��s���5?y������$���/ѡ�V�LԨss���E�"]��y�^����~������������GY`�`�_ta���F���K3��h���!")�l�,W�m3g�!�b��XY?Hubf��eky�Oa��r���_0'ٙ�iHZ�F+@2#�֋�(�
���2-`��O�9T6,(� �uʗ�*��b	��k��S�$��a�p�>��}�4Ǔ�:�NG�|�W^+^�_w+0sfA�p�����܍��l9P�	�1���Nz��7�%����X�^̃}�7G�v��#�x��R�>�GbH\4fG��'e��[�����K���疥R\�P[`+�T�����+ۜ��_g�S��b�w]�d�m]�+/3�[�B��* B����y���E|���aei�bx�v��gq��w{�z�3��q�ͯ�kw�n��ۥ<�|п�u����'�bߙ�b�xG����W����6�0ʬ�0X�;�7IWtQ�$֐���	�� �a[�Wa�{��a�|�9�<��૮���%(�����U�#�����o�gQ�����9�8�w����.�O�Zx_�0}k��B(���DZF)��W�\,3�P�������;;W��v�NqM��������£�2bxp�;�P�K{��>��wn��/&M�`��O:����u�(�=���)�ax���y�f�^xC�H$!�-6�0���q�M )���F����^�BM��]� �_��5��q+m�#T�0��z�~����eX>�×�hA
�����gw��ԀHh�q1�#@�G��n�����L��,�". �6؈Na�ORrѱ�A�er���p�����t����  W��8�El�:�A�=[��}:c�6	]>��e���iX�����D8�5�U��/��R)K+L��5D��#�u���{�C���G�-I��gͶ�3?�vc2�i1!�^Xb����~���*�R`6�3�Xd̯�7�, ǝQ\�LX��������gl��M��sUNf�?	%s!�ʎٕD0�cDXۉ ��Q�D��$�,��!�K��,��>̲��mN�$|U�ܣZ����{�s��P�xm�1�xm��cD5�餳�]9�}���u=��hUA��wI����҆羣����N��"�.�${�K��x-X���tϴ�,2I�a��U{��ޏ��yI���8�M�`��M*���m����j����^���A��*�]h ��g���q��r���ΗV�YH��-��?V���t�O�}��\e����8X�e�쉼ɭ�b|M��zm��=�,���Wα���ᢱ�U�tېh�$���Ό�qݢ�����E4�2q��?�Zk>u{A>��pz��kw��-��!$�H�������v� �~p!}�jO�OP2DGp2�+�a����)0���s�Z3�X�^����r�OP�Ni�	�$I� ��|����DLC�݋���<�������� �J}�h�ߖ˟}�5�-M�e;cyAhӦ۷�$8�����I��M/����1yŭ�1�"L�d9�淘��h�BbB�!�D�xYJ�yŧ���v���#��+����N:�m��ضm;�ضm۶�c۶ub��߿���ϻ�f�]�VU�9יs�v'����ˡ��kW�Q���V&�57�;�'�,�Q<��Ϗ�틿c{z[��d7�El�D������#F6Gla!�.gf_�)��#؋@���fBO�P��kA��h����^/2�p�h}.j����W��l��K.Q���-p�|���H�wMǚ��$�;{���W����5��q�(O�6#�/J8�KA�`ܮ7D
v��߿�Vc4n6�Z����_�#�a����[�(�5�!�TǷ,\&s4*�͚�j�����w�D<\��XX��N�j��(8jj��*�����ɦ<�}��歇c��2�`@�r���i:��F�
���l�v���#[�KYX��2��,��}啙��:��@��^���3���]��q�����C�wϥJ�͖��1�Ckɯգ�c{�<��)���~�Gޟ	�Ė�a}���v.�6��#�ŭbN�݊ �j�ז�*�"2<����|UB�E�Z����>B������l��Ly�E���gô�1�7YN�j�Kbpj�"[��.��,�l�� ������(���jj�O�S�e���u^�KY�.U��lb��6�r��nc6l�J�E��|e��Ygޘz�g6���o
��Z�����A9��R(}E}�-��@����zG�J�J�1)�T=r�*�]ln���&u�E���2l�Z���W���Z�b��t3�?�_z�72|�x��K#��6Z�+�@ĕB%�ج.?]RQȇ�?����#�6^sAƀ�>:u����+#�G��\]H�t �W^h�9I@���e{��; fW܎����<���Mpj������J�@g�-�,��&�2?��?�&��s��f���NW|ۑ�'�:c�@~���K�.�lBD���X�H��o�L:ٺV!5�#!�h�k�J˳��tE5.-a#�Vk�x`#A�fO:Dg��Ђ�W���,��hh��U�*!P)��5�]]��ː9��:Zd��ipSczm�����Յ���ӁT��'��a
ɟkc�Yl��k^L�Jm% ���sJ����F�\��_t=��f��ؗt�j	��Fe5?rSo��3��-��a�<�Vit�������'[מ�/�b����aH�6���p�gӕ�!Ӣ9낫L)��5�>�WPp2�ܝ�D[���G�:��Hu��/R��	5�t����]��M1k��RH�zbg%��z��j�2������&�ί�����[C�j  G՘;��ʨ���|N�$�m��ܲ��ư��:��%f �/����S��e�&4�����E��QP�U(�'^�d~��Ϋ??���#�tޱ��]�\��N4�X��H�/.����¾�(���d$���=��~~{����sʘP�����oA����W�z�i�
t6��~���y��1��*~ҫ���/��dv��.d���q��2��n��*%ܛ��Ӭ����Y5����^{?S���9'�fKu1�A��A��Q㮬�yGG���#���C͟�|���5��їoW����D��!*jW��t�i���}.6�w�L{v-�����ｯ��^�����8 ,Dq�Åɧͺ|��J�������d��;�`/��R�D[B\4����(ҩ%	�K���sH?c���Ң��~m�CG��H��*,���V'�\��k�<Rc�7��/�WbҒ�R�tO2��U���w��r��@�:.��H�/�G���6)弃j�D��X��	�P��}j��OaaRh!o(�x9Ҥ��H��A9��`1;�^;Q�6���쮖@X��aύ�3�>S�����������㛝�?%|b�o���<�~>\�1L�����W2�;�=��t5?�%�����g��U���{�f�^��Cv�ˮYH�n��$ݧ�&��0�S4Y�<N��ΘM�P���#jA� �������c�9�;�C��B�����<H�J�p��r{�3��x�\ҽ�G�!@`��T	\3SǗ��X���23��f�����gL�2�1����z{7#?����P��d{^���G����Ku�ϵ|�pw슻_��O�T*�f��p���سys�.��^��RF*��� ߕ�����#�<�P�h[�}�}Ƨ�8a�W���2�����)܍��5��g�w
+ˇƄ�e�U}NИ;<�T��BC�z٩��9�� ���k��.�����9��K������Nͭ���`4��qqa]���"S�+��:���B��έ�u�	ѥ9��+��J���υ���6(��0�^ΉZO���`��_�Ñ��%e�5u���=��B�^V��Z}}�n�jO6x�PY��^�����\�.�@3���i��uG���6��[b1��p�M��i/��JOp�+o�0�޾��~`� �Gvo�O�A*ΟW�#gmNs�d�̮:�,��*t
��'�����F�.E�VH���m9�G>I���˴��	�9ݑs�k����5�����~/�"��b���+&���\$�x�6$z��-�ZRR҇{ Br�B�;{yw��fG*7L��6���e)x�W>Z�曆pQB��M�`4&�}��Xbf��� l.��]�W�Y��n�}���@u!�S{�>3ƽ�ק��͵ڤ�3~q����^6��ED�E���L�k��~8��M�W�Ī���g��IܰRĺ^�уK�2��W*�����_�]�?\5�IN���D�u�.	oZb�z���~��?��P���EUg�#� K~ZP�U��Rl+hX画^w�/I]��By�fEƷ|�3�F4	��;K*YbVG�� �>�R�bh�=��;[h	W!+��v��9��G���Q9';�T�2z6��C��<�5C���zT��K�ܷ���D���-P���e��A9�l���e��J#��Iɡ����2D�����[,�����?îU$����HH6��#�a�������]CHA���|��a��ߵ.������׌��n)̾���{~tc���e�\�f<�����6S�/�d��et��5J��@�}�؜D�k.T<�a.�6�8I��<�q9"���������2��GCM͌�nȮLƭsd>��:���)��C�J�	��Ńڥ�~N��
��qIQ=��R��	�|>��cم�҃���_��c�����ʹ�Kutc�v�	������0xY����@=ד���� a�b�9�F�K,�p$�W	%�QG�;q7i�(Si��� ��s]2 L������x�[�_�5�ح�h3�BA�.�R��T�h��!�$�-;gpڂ�n�1䋠=�z����~=��@��k�ջل_�٪�F��c�!c��r����Wu�fD�}����P���*G@�M�L��ߒ;�D�:_���~���w��yh��_�U����0�9�,)gr�HR$��H�L���7��"d�+%�_pl)Œ�5I|��xr�abF~ 4�э�A ��9�⚨0���÷��f��,y���|�;��L�lt.P����b]Rpgͣa�}�;��ϰef�Q SA�<(�	��K�s��]�ߩ���nh6r��K��:�3V�F%���)ksB�l�6�9�@�EB�! �np�_�[	�$�7 U�s��_�)��͸=:�K��)��_RK���<gjf���a��&�cA�?lЉgx ;9q˅��&�JQ~[�ļZP�����9�}2�����hW�o���?��u�sLM��B�S(��`���[��f�wr�H��`�;�(o�x�����A����na�O��u�KM���5CG��f�*)�u<�N����U�J�~C��t5Q�Z�C��CH6!G�͂�V�Eѐ		}s&	�-��*��QX�����T����g�a�sc?���)�;|*�@�Qv��h�c>����}۱ ��rzB<�l�;��G��������K��i�.g�Iu
���ة��T�?*׷?����SB��Hv�?�'���By�7���V0T8��׶�}&��#n�n.\d�]�����0����n� -w�I(�%[�Z�j$et���&+�^���L��0	�G$�{�+Δ*��NX.-�v�U�ޚ-~k;��c�kmN����'Wu?#,�Us��*Q:�J
�0�"Z�yE�8l|R2���S��bZy%�
���Ke!���pRZђ�S��WB�1,��4�hߕ�VH���(�`Q��a��Џ-�
"���P
�/����Ð[1�� Mdlwʑ��'����د.aE����PG4�,�uĥY��O�9!�/Y����p�
���Z���Ufr%$O��L�RL��"��ߞ8U����}3R�����G�뜨�����$bL�����)��#�_�"t/(�Q���/m�A!�]cPã�f���T�f,*7m�3t��2U��D����I��<􍿇#�E�ד9'��2��#d�+��X��������Na�g�������� �ErPE�O/[:k~DR��4��F(՚߾���{�B���j������O�xopy|V罩��4�索^Y0z�}�wQ/��~����ܫ֢SNJ7ن]n�11j�L�J��ˋ<�K���
o�ê����rK:�j�;�j���iј5/���?	`m
��Ȃuk�2��ۥ�����)�]M-H�i����_���K{L��So����z��������W�)�I�~��Q�z$OVF��n��\=���yvnƽ�-�:W�u.��Y4�y���R�ɲ��x�8��"oB�Fػ�%,�*�E��??-!3��RdK��,�:�6�;K��l/_8]#��Ã�}�.f���Kk8붃-v��|���9�W�KNF>�k�L�<�I�͖E3T˷J%��?�(q�#uh9֡�ى��Lg�|]Ko~B,�1��0ֲ;w�U�bu���G/2+�J���T�m�Y�6E�(�+�@(�U��yi��@I���n��e(��]Q��RL��_�b�hn�7Ew�a*5/}���9���nE�ՓN����V�6�67����G�ݣkN^�.{�Ā�Ҕ�h��9�.�T7����_��y�u;ҍ�b��P��BrD�z�.b����J�狖͆J�>���Y(�����:��^$�]*o��*@�)hwzϪ��{W��q����IQ�vDЈ�*s�	Vb�T�#�?��}2vd/�Ϭ�c�ZM����:�n@=��R��3$F��^���>G[���ס�l��f<ŠK��˪6��6k(��F~��.�`�h@d���2I{�e�LĵXr����:��Y�j�G�-�,�zyz��d��=��]B`&��A��ډ��j���q�K%uT6m����z�+e�m5�id���9(��)�V2�M�aR�*1"����x<�C9	C�/uz2��[�9��D�9F����Po�)}��S���Wο91C�mz�:=�v�ipS��r5��Z�l/�`]>�N12�ةW˟ݮ�}Fu�u9���4^�I���gg��TM�ή��?�Zad�Űa����X-Ew���ydJ�d�(����+��<��g�x�u�X���"V�B��Ki��C�+֞��c��9�l'�wn%+au���|����	 4v���c��Y�:�f�/u:����.�\��N:�'��h�Y�Y=�&�Z\Njrq���׼�V��7���II?2�)�B���M�-�:MD����Vm��S���J��4������/������v(��Z��v�=�<���ʵ�)ҵ�$43n�Q�t}b��##�B4^"F&I(�!��[_�)��:�Sx�!uU�a�u��"�m˼���*k![�dH�`�g!�n�
�+v�4��o�b�7+G�#���*�\8I�/G3����#��
�77Eg7�����Љ8c8�<�17)W+���Ԝ��	;���ߠr!�Hw?��D��.-l)�,"c�%M�`���˰Ռ>H�v����r{��뭁�+�2���>� �i��u���#"R��/ߞN\9k����y(Ҩ�`i��9���6c)��qF �)�a^����9����gBE	)m�
��i�o@$�--��l9r��q���No�t�B�}b�B���G��{�15���+�-�CE��ܹ������4��T�:����ݼ�'���
�.2���VECu9��M#Ak�yC}��}�go����^nU�r
�9��Tv6'ND�'C!f�w|�n&�L����!�&���8a(�h-}`�^�"�eT�n�o�5f�j@"��-�D)�'~pz��`]�T:q�gLň&�]�f�j�9Q�`L�[�@��n�Ɛ�)��aS-�l^E/�����IqyFy��z�	��I�Hq����ex�%��������~�Npr�fǼ� �Ip��&a-ʫ��Hd�����RP���R��(G�4�e�^7`a+,�F̾�&��5�{�R�?{�pَE�����kR50U?��6�0G�r~)����*����G��9iq����_Q�Ub-'2fW�h��]}��]������x�3	�w��e@}W�����ޚ������X�y���Z���$@lL� �R��$�Y[��E.@��
��H��GL��y��_E������tJ2�o�N���uFf�I1|�g�dZ);�Ģl&�̠��V+`H�N�|qx�)X��^=K�U�.��ˌ�����Y�<7����}�1sLOc��;J�
��vO���J��4�O�A#��&�,�ê#lE���E�O��W�X���N�Δ7��Ԉ�.�L����eh'�d�f��k��o�������+����Y:y['��j�9��c���W4o���ڽ��᲍��t�l+ h.��!�,�Շ�߸̛��¦?b�$��$��&�fe+<�z֧�/NH�{�(aB��ˬ�	�!�6)�IE��0�����<ax��^����I�m�쀫J
/15&"Rvj�&�\���674�i�zsi��_+��V��������H%��MA����KK��A�p�0K��p�@Q�Q
F[H_.������XBK3�����ك����d���K��8:���A����L�C��Q�@�**:� Qp2��9��4q	�:�*�d c�0ĀX��4��U�k'2z.%��0��{�ܞ�et�� �4���B������,ʥ��e��ZJڣ�{#V[|�3���?a(hw�tDA����a��er�k�}��$��KrBK��5	o��� �F�۩��<��?όxD�Ϝ	E�\�4+I�9��L+XsBa��l@�?|�
<"��@�h�V i'k�Ü\�q�%��
�j����7��$���H"��%I+�0�5��BY�!h��O�M>$��'����ܚ����.� �~	���h�PL]u������ٯ��X.������O<fX�%=->��bE| ��z�P�6�}=`��K���z �yѭ�;xȠE�t�v���6�����8����o�I1�|��8�ޭ3 ������6f���3��F`�uo�=��ÒfB���O]ݏ~2;`�f-v[2����֊�����)�f�{��S�t�������3�"�(��a��1�b��G��	�g�nX��H�P�X#�Η$���F��Ӗ)*� ��5�ʌ4�����r���Ɓ����~`c$$�0_o���缰A)���a����b7������Д�_Uƙ_:̔�����|� �>S
:�q�{$#���U$��#~AE��}MF��X=~eIz�7rk�`�����z-.o���?\��_#E�Y���څ���;����Iý������� �^)��*y������'W�����q�@�����on��@�-N�se�U߲�+��F/���m����}�NEV��'1��ai��N]��:6�+FN��7�9h� ؝W4Rcd�����J��D\���0�����T�Yy廎_�ߨ��dP;���-�&� �u� �F�����hԪ��i�E#O���'�s�pPZv���\��@ƅC�l�C4��7��Mrk$�)�c��-�
��6)Kt�u:�E�s�~�Se(M�k��X�%��pX�d���\�
�M�|�f V8�"!�����8��/l���)�;���o�����~�]��ghlV9ƝG'���P�L��+�ƭ�,�3�\�8���~3�'�[�Tݠ�N�q�rLp��ֻnLO����m�~19�Ģ��&_n��������-�w�&q*s1����eׁ���`�I
���N��Rc�.-q�����D���p�:����E�l�bڣ�󤴅t�+�!R�/Yf^
�]Z�d����ā���]�e�S�w�K39�H�PsLz'
�X�g��X��� �k�쐷��q�h�Xlݠ����~��J�6���sF�$��&��K����2h��J[�\o�W������kD$�)R}F	�/]�̈́b�B�hA��@���y%\ �aې���TŖ�|ܘ��w���!\�æ��A���Ĉ=��}���׏$��h�|!��T���_�� 	M�1���'d���g��aP���5K^4�����(������B���!ne*���T�Mv���&Zxlƞ�m�,إ���O��As�O��/H��lǿʑd�L� �s<��C%�gl.�o�gg�$��{�ܹH��h/a���I���\1�)�x���i콈�D����Q������6�?|H*d5�]�R���¯�f��w�4�Х�{��"��'o9���E���}@Ү+yL��J��>�r�����_�[8[y�����th>��]�+�^loM��R��}����z|�)m�pE����(��*�,��uS��/'���sfq��S�-��,.����!�U�p�E
1���.�_%1�2_����2p#��p�����k����Z*����E�o%�b�L�Rf�,Wпقcw���\����!�B	�
(�'�` ������6h67\Z
�������*{��2���t�e���u��ܷl��K�\h��ց}�H���	Qñ�Ƅ�l��	5)�њ�[`��U��E�����'���q��
L�J˭�P�O��J�C���)�)�����U \���	*��ep��S���� *L�y���.y�J���K0��Z(����	\�F�=�G�E%@y����qD�vd�����a��Mϔ�ȃl�7X,Kɻ?G�t����r�p���� �g,M�;i��?n����탼�h^��8��9�h�4YY �x��|��"nPPPb6B!k%�*A��,�z�I�E�\+�HO@��&$�<����G}����E	��ֱ�~�� �_ګc��FL���Ӯ��|���y��,ɭ�����%NV6y�@ŋ���K�@N7(�}u�\p�V<��XZ�竰����l��E��9N�A�������gl�gn�p
�'�V��+Ж=)e
�xDe��_ug&iG1{�����Q�
�4���]C���q��Xt�~�� �G�<Rք���M���X�@9��		9��I��w�N�s�D�e4I6łOy	Xp�w����.�W�|fr�?>����/�����W��3�[���l=ͨ�]-嵓U��-�m��m����t�&�.��i�7������GRk>����� ����Բ���bMd��J*�q�V�ʈ��ߌ����O:����k��\��_��q 1���q? �6�g	��R�� ��xQ���Y5>�n6��xnW��x��wר���s�E9���<���I�)<l����ϷB��Gt��0�B\٣��-:�i����o�,4HR5ॱ6C�J\���٧��*nUT��I]T�'���aO��
�/DDL>3�#��N@ٸv�eMq��d�c�����;���VC����ˇ�+���#�u�� uVBh��.�T�����b�h�����>�ж �	���⻮C�6�fǉӔ����3�t��z�v(8��xD�<�pf�{��<,�$�u�Î%���'T݄��sKQ���@��8��l4�)\I��J�.��h�*o<�hkNdZ�X�@��-CXp�-}[DHW��nҀ�L�[�4�`tB5�I�<7�7�)}�J�PKŠ! b���)��L:��h!��ͥ�l��&w�ǨK.�V����+���;8,�~�s�g�"�Q���ۊ����&OBx���^�^_��e� �AC�NЃ�꿤a�"D�-��.��z�c��<aˢM�]��N�fY��?�!�G(Cȏ��p��;�m��'P�[��0���J�f|Ӡ��ƦR�Ǣ$���G?s`0&�4�~dg�ļKي���U+"������$fpH��o�0���`��mN�*�.;��f7}�J?�.s��A���B̟4�E���]v�q����ĐVm[Zu(5�<ic��wnq��yԱ5Bհ��o1�����P�*�@���7 ��V��#)���	�	�����������*-O���ZN��S&��X�ۗ0�U:;����n�,B�]&e�	��1�8'��s%�Lt��.?~���ԞV��夸0��:���J���@�q�Rĥ�B�����."51��N:%&�y���?o�!���xF�k����V�Y���BֈB��S2j����kE������@"�`��� -'��]l�-|���r/I��3���y��j�)�49*�n���1���Ȋe5�-+K��c"L�S+��Q_N�onx�0�6�:=�I	�YIr@[�`2B=��/,v?	&)���s
��n$�I7�;��|#��h"��S#bil�-;���N��S�	���<��}�'K�>p	��O_<	�����ƈ�w�P�a�����r����mЬ���ȋ����g��g��&�*lo�^##�A3�SY��-^�,I(�3�ϛ6�ue8���
@G&�ҥ���k�Ȩ���i�u;:������N��I�������m�L��p���	p���x�2�zh�ܯ��!�sM&��` B#zA�B�xvީ�-��a;���j�h�*@�i�'b���9��^#+�q'+��Ǔ�D��f�z����}}$�"�9�P���-�hSB
s�H���}@�R<&��:�D�ĸ$ں\�N{l2�&��B�u}�a3~R��Mk��B#��	'�?�Ys��[q�B�W�u���F9���I*��R�P9����p���Pv��ݛn��l����0Yd�+l�[��99x�򚝅���w&���ҏ�ͮ]��Um
	]<�����`_�V�*�k��sRǜ�9�}>�y�ᇆ����Ι�W6j�5���.I7�v�����q�×L�);�Sa簯�D�iO��^�PhW��ǥ�Q�u*��}Y���U���#ο�;C��*���yp�swJM�:MeWS躜-q�t;�H}���=t�͊-þ���h:��� ��a,lΪ�)��mwV��5f�����Y\�+q>�0
~G����Y%�M��B�"Ū�$$l���Q�g�X��VC����ߚr�AF�|X���A-{�� �*@L��/��iM���f�E�h�u�����E��d?��7�Q��� �2<��.t��3�i2��?	q5|�PU���tIaM.��@�Eu}|��9l��N0���w:� +*Q�	���V��H�'��%�g,�.y��⣅��}+X7x?���^f���Oo���O?��>���_��ۻѴC���E�#ؑY��i��g�:i��l�XF(BR���Z0d�e�W�.a��=F���q�l�z���A�P��p����������r���Q&|��Qv���R3�b��Zޑ5"���F,�I�chc���Ԕl�z-V�(�؄����������!3�yq�T\8�cMV��U����T��x�2�v}��{rY\ZX�*�S��I�\��Ѵ`���,P~�t�΂V>��1g`j�����^�'���O���y��Ǜ��<�E����BY�K�L|���ǡ\wF�G��u-k��h5.��	qg2���h�����Q��`�s��ڊ׏o�a@���S1���Ÿ���.a��+ t� F��E;]w���������qu_ѦL��|�HK��{�K�]��#�fgU�&���x5#�c���T�@���2��I�����@�ϥ�y���X��Ӽ�n0���T�{�˸�c�xњ�S�O^�O�h}�{؜d�N�週�nV�\��wPd��?�$�8.����|��ޥ���������D�_�8����1���L�f�@ǋ��i��Ճ���`Ej�bꡇ�"]&����>�S�p�k�96D-d����ș��V��L�]�6��"Y#�پ;�:SN@[���������٪��ţJ#\�t���&7q���X��B�@t'�ۺ��3[��<�\���m{������j�ovx���ؘ\_�0�5B�:��^��>U(���U|-�ӭ�"��F����6�W7��l�����4���_��������K�	��-���ūD5sl�FY��ߙ���������],����Ʀ̜:�n���'#��g�J�!8�j}�I�TZ%�#���ɡ�)n������!����t�a��F���LuN��Q«N"�i��>��T#�ny�RO|{:u�%��L�|w�>{�6|��o)���L)4���.���9�z�	P�}�������w��~���Q�ײ_b[�� C���%�d&���'թݻ͈�Р���X�]����c��`�r��9ί�WR�7�j�I���I5v�ח"�b+2�����$F	����é6��epa U�3��	��J��'��bt'<$Ǖ�>�c�*h�5b>6�sVfF�P>/U�_�f&��ܶ��S�����X%���'��Ib�C��݇^�+���6DD�_����tW+��b|��Z�H�[xU���em�`��UدI���|@	�T�&Ye�4F4�
�#mE8�M�i2BrOQ0g�^a��:g^iA����]�M�� Ny�	�\�_�\1T��o�T��z�k1�=���U�&�,̘�H�G~H�<��ߺ�祱Yv?_��Q�����i��=���T�^;��E�|� ��5�Fc�O	$*DU={O���ݷ\�7�ա����n�[D��B�z���x�g�b�1�s���
�B���	���K]q��Ib��1"����(.��zE��7����U�/���o����-,%́�dF���>�i�iR\�CG�+;m�ԛ����{�[�	@V@ 6�1���IT|]���O�K�@�M��	�=[�=�[g�qBbl�>�B0+�'d!������СZ��vxc�����,��5	��������Tb�V�E����OG	]N
� ��:o�U�"ާ?d���S���\?�uݖ#dG�
*�t~���ޓf�"��F5"�p`[���T`���L�J7�Sqw����b����sG�D�|��<+�P�F*����9�nP��D/f.y�rVI��a��!!}Z�y��#i�.5bﾮ>��j��6~sHLB��hk-X�̱���K��Ml�������I�^d��1���w��˥լ\}+M��幪��K����S���p8����p�����bR<xHB@p�\g�U��D�bZ�
��- �bI~�u�V˸���JuPh�-��D��� k5U#�\��~�f'S��d�"2桽,�¹w�;_F��ͷ�-��0��C,�5#�������Pa�H�RVÏ�5�?ן^2���Z�%K`�g���Sg$���c�I�Yb�1b<$��Ɍ	�'���廨߀UR��2��@�@`Fp;��$(��i,��G���x�v��{����!��P�h��9dy������`L�ؑ?��t�ۍ�Y�]~R��
,���7�h�&�%�F]#����4R���c���5>8�yJ�=g�d�D�iPH�\��FuD-���H���N��4x���4���l5��h���a�W{mY`	�R�� ��8|���%!,��+�(\u�k��h���.
Pp�":1c�Ky�wYx,�yjt،�m&v3rR�hӊt�^D@ŉټ��E�Y��'��G�\ �(xKN�.�����8������������iO����`w��5��'<h���wm���AZj���_��3��#���׻\=SX&|��t�e^�#f�5�S�p�0,j!Twu�\�0l�mx����;Z�_�6<���B]A�ʖ4�U���Ebd�Ь�g:`:r����s�|�}����|1��D�G� U'�TSƑ����@2&% ����h&T4f�?���k��hO*�-�"N<8�;d�퓜#�H�Q���xf��]Z��Z�π�#���7)����}�}��X����z� 1B�&��[F�|yf���'j��KV�zK ���Y�I�4%<��8b��PN~Y�p���AMi:�p���(y��4Rm�����h�2�6�Ĩ-D�`5P�<v�I��+�������ScB����%�1fV7�m���22I�ڙq��0�#܆I؄o"M���>��Ѱ,��b��	��7�:��TF���&�K�?�'`��Ϛ�RB<���$��T&����%2���WD��W�cjPg���+(��h��j>�}�i�T��L�p�pi8k\�=g�fǥs|��9��	y���k}%�+~4�L���E&FkN�<Sp��Ⲁkŀ��X�6�[1=k�"��ت-���I�M�4jX�H��Z�F���ly$�Z}s������&��!�C������͒�yS���fA(�	~g0抑wXh�Cơ)C�P�}"�L��Dm�)nŎ�.��] �l�&�m�ZXzЬT�����)�f�j�ns��H�����rl�9oyޔ|N���Cl�n4�9ϲ�d�Xy�T�l\��qTӀ �F�9��n*=��	�7��iV�1�W�'b\h�D��E�p��)CT�=�`�EUbap��z;�6�F0
���@���� U��se�<��PND�`hL� jJ`$�2i#�b�@�3�?�q|�2!�$[������X�"II��\}i�<ʮ�^?����G~m�>�������F����'z3�͂�/B��6L:y��'
�12%@5%y���/�d�%�f�"tZ�4�q�V[��@��KKݴ�t��T��� c�m(�MZM<>��7>���)��r���c�Z�

�+�?J]xG�Tf��YCp��l��x^��цE$�-w��m�q-�I�G�����,�D�M=)��@3��I��^�QS��|�۱�*��,Ӽ�8Eg��]6�G�c�� ��eÒ�ue�_��I���TbO�B��б�i�,CP�x���J��<$ ��,�l�=7{�w��	���`�5��H��W�z�_j��x��.���)JxI$N�Mͯ�hn񲣄�')��J���d��*7�q)���XKC�����d�J^������1��ٯ1�|��n���P���L���6a���4$�\�&�q|Rvg���p� �4W���٨��d��gd�#G�yh�����&��3�w�ї�q�MBWy��(���D���O�'��O�B������1g��f&>Gq{�X,]^;,9�A����G��lj��0�Ɲ�,F��8&WiQ5�ٙ��*����j���	Hh	[u5!�#e�i�U*�^���ů1_oN�exD'�#n�c]�po����J$�.�Q���?���b
��4�]ơI��ɭ����KͲ[0��1l��-��`	;G@�#�;B4�ò<U�����F'�儞�Ql�;�Ѷ4G��&/��u�p�6xG�H�q��r�W���w�?�br��|���1knoˮ�?�@��8���Dr����f|b��Y9e�Q�ӡwӉ�@MV<
1�=/@�!��"x?����?��Ȏ�S�+&�.|�B�Mw�E �d�vS��!�mW�= �{f���î�$o*B{F�\�	~	8Ȳ�Ԅ���F��H'-�,�B�M>�e���߉�"P �tַ`�����tC����іjM�LU�-S�f����E��c�<KiT�yj�g��3�2�F6�:U���s�f�3 ��X&�v�stMN���)�h�>D�X���qɈ��%��O�y��2�Zr|^6˰��$ؓ�Gw4W�m��.�,���d�<*��g'�o������!c7ɮ0Zg����dpE�m�w�,wI������؀I�acmxW��&�H2�P��	H4�gF�y��� �)|��b��ޛ�M��X..���ZR�s�=� e���xJ���'��8 iB��˗�5��A�X����[��b'�F��VM;���u`=��wH$qBBHBB�8~��������G�U���4������-8,��n��K��_�5�k� ��;\������:S}��<U[C]^+)��)��y6����'S՞^g�y��=��g	縓m�����h_�-H֏ �p0�3%3�z��o(ӕ�v�̳��]#N����}z-�@�hi><��r��/����e�R���gΥ�z�~ac��:l~-	�f��{����0`$��=!6�؂nOĉ�B��	��*�Cv�k�u�KARx�f=��Q!�`�/���c!ƞ��q�$^�x���ኈ N�%��/a�﫭:�ϕ|䧢�����JJ�P}x�P�|K0��M?�.è�
M�������,%���u�W�3�����ø=q��A{�_$���$����&�:��q��3eŜ#�� Xm}e��w	�iRQ��Z�� ��@����Rl@	���+�U^>��%.g����p�В�B�υ�0OO����OOV��D���E]�X!�YIG������%���U�	�(����B�=������;Z}���}Ǎ��T�
l4�y�vNM��戺|�L+$��_��:2��~�#8.�񁩾�����b"����|N�-�wX�\�a���f�e��E�52P).��\��M�Tr�O\�`�z���?�+A��#^�~�Րױ��ng�?>a?i�����C��������B���.L����[�����m��ը�V�M9=�!����]��iX�8s��V��>y�}��
�<Sɾ!�y�p�1�IB���|�M��B)��<��a�{���v+#���7�jl'�8������W��������������3�n�g�����zs>���(g���6^P��e:u@��/��M��a��w\���-�.�Y�r����o��$*3�RՒ�'HBB֝X.V+c���k��=�r�Q�dw�Do���ͭ���;E�,��7��Q��ͥP�4`lQ��k�<�^�ɬid�T��ktuW��ʅ(�+Z�.���d��E�Pӛ� nDb�TG�8=:9u��~�)�ڵ�Cg��z%�8����P�zsf~�z����D��9�Րc��&���	OD���ms�WvC��P����������W�]2�s$��Iv���ͤ�e]�@�~�i�P�݄LI)�9Nu��@�h������K�Iq���Kg��^�FV�k8���"b���u�^�3Bո��.��Yح�{��>{EBh�g����P��5���2/e����Ǝ���/�Q����0�R�m��	�ߥR�.RR}�	k�L+EJ��:�������:KC�I�W�m8z3��n���ˆ�[L��pMH�\d�PI�+��d����C+kѷ�9��ݡ�<j��贍��:qWF�d���U�0֒0cR��?;O���^��қ��7��Z��:ێ��{�B)��31Z�m�N:A���˛{��*oa/h�H2Zo"��kH�4�//��j>���Z˙S�]�F0���ղJ�룺<+&����T+�uC/%�7�.���\TbL��`=�5�n�@�ZW,͍����$ 	��;����H�!��<�e��(�[
e��5mg����F��D���v��FI�����0��"��Yi�sF�ҜD�l������^ȾM �l��w,*��>�$p�F���2�����pO��S�x��GL�ק�/X:N��D�����u�h���)Μd���hxd+�t�1�|����iil�L!�dT����aav����THv��	*[���x�Æ�so����f��8�l{��dl99���������������0����{�?��EN��},�>X�Q&�O�ID�Z�aa�P����<�����A+���%ѡ��� ��(}�i��z�y�Qq���[+���&������������V�]U��滵��?���8��F(�� \�L b�=0@�@��7��쫐�E����|��n�2:�)�����cW!�'_ty(��w'B�2Wv�_"[��B��ZF�/��&�-���F`|�L���9�@��#��Q{�0����6'��OLӨ�eYe-{kr��a�V���A��p`Z}�����aOqGD|�s̞�Ƚ0���q�e&;��m���oҲ��|�����|�$:o_�,
�;��Z�"8��r��U�>�0�������8��1ެu>ry�'#��\�j�۞����ú�gg�V�h����Z���J�0Z�XwR���^������7tW��R��2�����Y�=b�K?!� ��zQ'��z���uj����6�r-ǐy�"�(��CV�8�4����Y�3-��^r���Y��ab��J.�S( 4�Rl\\��G�fՏ���%���ʃ{�>[ ����ujzK���w~W�F��=f�J���ΥF��/�I�9�����b�4�UP��J�^`^�=� �u�\�;�볕Rl�g�l_���(�������M��^�f���?�c�<|	4G�s�X�O$�=�۟<M	��y�"��	�Y;��\�h�T�Ud�3�'-e�l��;/
 ��c�Tdk�"�o�;o�f�'JA�����Z��;ę_��p�تD�H��7��:-B?}8TJ�(&QZ8P9B�3��&q;Z�˞7V�v��0����BI�M�.���k'!�r�\N&tk���R����Xv��m������h����>��J��4$��g�����f;�Xy��"^�ޅj�ּ��!��NQ�Xm�Ĝ5���!%&;��cPT�N3ieX;�`�xw?޵ ��yނ�����`���!D�-G�v[�bR��HGf�����T��N�[W8�l�>ѾY3f��0�2����!q�7}�!<��g��AÈZ�"�����2\�Y�����L�PÄ<�]uB�L�!���_O�C=�˱�z�H��7�.k��h%��ާ2���k�OF«����y�ҕ��Ӄ���}@�u�8�V���*�魨Q{%�=�E1�@��M�ڀ̬Ԉ�C���柋-"ۂ�1���=�Y���;�=�8�~}��ܽ�h��;-gy��������[o�g�C��z��>�.�5��� "b�|~*M��i��!�+�<��`
 ���^&��έt�\ꝩ���B���O�wU5�N5���g���-j#��4�����L^���t7˛�7:7kB28�z���ۗ�Z\�3 !�i�cd�:����\l�h�\�4����U����ꀹ��F�W�sW>���}C���b~�J.�W;5*eQ���������{��w`��Wt �g���y]�R��r>^�r�&�t�)݊kO��~�с�����='ov�c�v��絰����k����t��K�P����gr��,�)O��8��,zjG���}��j9VM�S�w̺�������PM�ޕ�m�G��(�_�������?�֑Sf-'���rx����*����x�!G �1|���b/,s��F�K]��͊R��tX=g�*�y��ʂ�����>�%ǝ��
P��XfU���Qs�����y��̑�۔�7�����vJ ���l�&k�+����u3rƔ�>a�����!���Gƶ.-�Tt}9U]"�� {��֌�&r:]�����l�ɔ�[��Ќ5��tDߧk+��_�~�cR�>��;9U��+����a����&b��c@���~��m*��a����q��
`�X�f
�*�E��|�x�I&��j�jG� "��iǬ�@r`��{\%T�n�����Vk�_g�O_a*P0�N�[�[׎q`�[�@�XZ�1�cH��c���ڛ9i�>��PV?C0@���r��}	�I��Bo��*~͘Y�gtt��DS���	l�GwV1�π�?���Afhg$��ܶ;ǩK��K�s��A?f�����|�&��\�fۏ�)����n�R����1�Lx��c�@���Ɛ&ꬷlm�
58-��Wޡ�3t�Z�1:�N�']#:qt�X����ɼrMuSŬ@:�҃��EF�����h�t�]e� ��6���f0��%rY��'�\��!�uxv	��>�JL�:��h� ��9�t��u��B��Ck'����p�:�}����R��y=z�_���`̘���*���@�{NU��$���hoX�;��\'"E��#��~�K��k�h+�٪�����7r+F�~ ���"���4����� �1��h��K��M�cX^y�p�c�<@�@=���Dc����aot�4C $F��1N�L'B��>��؏�z9q��20=��ރ�����r�!�_�_6z�����sm-Р__~����"������u��� ������kG�i~��Fz�[��(A��^4�l>��f�>��f��TH�"H��~���'s5����$2I�*̓���/��fU���<BP�ep�X3��pEy+W6 k��/����KZD�n��9��b�3y����x��5�<���{ ݫ��_�^�ٯ�ٜ�Sۦ;Q
bȰo,�g���j�<@�p��q5>�����$�
$5#�[�+a�s'[�DP��z�b��%��K�k7a(�+��3���x�;�ư��A����`@)��� ��O �h���Q���' _&G1�n��G%�iD�&}�����*�A�*�jJ��ғ���5�����ð���^_'AB�>�X߫���ea)���^�������M�]����O��Tw�RWl*���I���F�a�uةl�.�h�<�&7�9	�
�C�8�q�Ns�	��l�u�u\aǦ�g@u)&?�"5�0����(�Q�� )	ek�@��T���&��J/<.i��,���^v.����-Ύ�o������v�?�xO�K������$c���Raa�y5?ck��ӝ�����ru�	F��Q���Mn���-u^��}OJ��yX�u�B�٦�yJ���y � B:���Y���/� L��t]�"�.��x��p��dھ%�WO���w�;5y�9	 w0w���b�ο��k�+3��Z��\5��z�b�N��K(�4��Q��O_=������d���q�5Pz��a<(3O������j:��t�D�gW8�dRnW��t�`b�rtZ�8���K�3a�u�y���ߣ_i[AX�P8Y@MN��e|���g����T� �䛲�l9jT�~��?����>��q{���}IǞ�J�g	�e�z=h��y������@0Ĕ������̓p1<�]@Ñ��2s� �#O%1�'EkO+��u�Rh��do��eRYl�ԭ׸2�xuo�I��q����W]�a��f/��_P5{�TpVœ��b�j���͖�`�Ig�OU9ݥLi}3�����wG5G�l�.՗츭p)�|i��C�"	ץ��Z~�p!���F����N8�#Ϸ?[2i�)��c���wh��rާ�d�(v�4\Je����J;��0���y�ϳL��%7�Ã��o��55I���k�(?�e�fb.�1W�G�EIHF��"�s����WU����H<s�X��~=�H)��G2n�6Y;_�]"�[2��h�'\��
sSax��ܭ2N.ZOۉ�~���������=>��Ы8�������]�x�H����iʽa�	�G$�jYS��8޾�]k~���d���o��Y�:,�W�$���ֻ��FqѴ���l�ԩ_T�x|�CI��(���7[���\��v��m{��7�P1*ћ%H2�=oSh.�_���#�ߏ�~�'۠6���ܕ�<��t��8j_���Vmu��%�t[��1��T�N��Z�䖝{�֛b:~�H&7F���a��?N-
TE�v&6.��� �x<���0��^�E0�/z#��}p��G�ArK�"s$���7~Ϝ�^JQ�>���֠F Wzʖ���dP��ʺR$h�꿩��%�����L�:���k�e~�&/��WO�گ;�~e�� 48���wQ;�v�#/�^�̨%}�婣�/݁��yI��@�y(m�נW�
f��XTZ'�@:�'�m�xc��C�Qq�#�Ӛ��3L�Ux�o$	��cB�CE���O��F�I�5(Z�����t�%�D�a�z2K���\uO8������(�����>���L�r̝W��3��O����'�e�\�o�z��*\"����DK@�a�)���lJz����N�;"��ǒ44]� 7H��T����l秫6�>chd�Q�s����#Q�{�比pD8�ԕCx(�K�T~��[q/�a}.�y�_��*����FL����F���Ŧ8~���
]���YPbTX�F�0���2rW���w~�B�Kb�rS=�>�~�Gw���ao�N������˘b�`��	�|�����7 �D�0� <?n���d�oR�/>�9ȞH��W.H�O���I3~���y�Y5 ��f��5S��	F�#�c�;���$����4~B�f���BQ"~y� "��\���E��__Ɨz��v��>���y���~E�T��b�S�i?����5M��N��˼Y�"�dۤ����絃�,c�ԣ �b
BHn��akй���df��������T����f+�!~<��G	Fi��7؁���Qͩ���oxX�Q�vJ� �,��� �>4M�a�ɱ~ܷ���py�U;9�St��c{ǩI���L�6�7���&C:��;w�zd􆰧�oQ�.ϝz��,�_��[���Lٙl'h_.���|P�S��65���W�fw_���u�y��]E������!�B��uH�2q�Pȱ��E�%ڮ@�&C���c{�������N��7���Sl�}�K��C�<�Gd}]~	���T#�_zR�%�_}���hl�T�K���}��n�}�"�����a��[����Y��u�WRd,l�D_;a�7�D���\��〭e�?�-[�=���W����l��m��Н�}#gܸ�t��~ib�o��%�F� R3h�}��;w""R"����2D�e¨������E|ҝ�!�!ɣ���F"������M��6٬&������+��E��.@�NåN��Õ6�u��yŢ� ,��&�|C��\�:3���~ZE����wR����7�?�#%�A�䠩mpl~�;�NwQ�m>T]S�_��q���h����������00�f#@�Y�'lGEA@0Rh�+4F��,VF?""�)����ۇ�>�0��ϼ��0q��u.l�w6\6�4��8rI�$%)y�J&ťN<;Z���ϭR�Ŀ��	�N�%� �&s��#��� �+*�G��3*��B��io�9���mX���f$^����g�C�5�6����Z�ٴ�, �Y�MC��H�^L�5'������l-!�C���8F��.�닎��FV�S@�2o���ߢp\��~	E��ўz`/�yV�}!����g?u]� �<_-}^���V�z�!���}?P��g`��W|��{������;I��!���Җ�)�㸊�������q�X*��U
#F�%��a�C�V�=�m�,�39�4��k'|#@���e£��V!^F�,�W�4���C�u+6�Tn"+�Jh����}�ؿ��O�:�l<%u�UÃPtwR����ÿ�T��;��5�iOx'��J��N���x�nB� ��Y��n��JF���vſg:�I�y5F���-�L �"Pw�"2�}?�|�u��e��Hj��Z�"O]h�����'� �&Uh�4o�E�Z^��jK�н���3��Ƿ��n�Mf` ����(�yi��W��td�q��ޘE������[��OA�U7��_�P���T�aY�Y7c�
�2�p�T��sz|����V����N|z���= ����i���c� �fc�&�W�.G@��ut�cwJh��޳��G�ʨ��d�����0��Y�	?u�Ơ��X��'h��5Ŀ~ސMDeAW�̡���hr�|Γ��Z_���lWe��B��MԿ}p��o��PP�	�0E8`�l�A�k��X�dM0�O��zi�������_�]�MҜN�0D�v?)AÜ�g�l��t�IW/t%�܀,���5��c�^rGafyh�e�bWK? �lf������x^�k�e��<w�-��Á&�ְ^[��p���w��\J橆��A�Ɓxy�jb$�f��yWnz���X��j��c�7�s���Lx�BƹC�R�@�R�����t�������W����KQ�G�=��9��$<�7"�<���n?����Y`{Z��v<J5g�ַ�i��Hu�(��I��Lq������=uui���N�b����۸wͩbS*2��N�}Z���#6|� /�U�н�m��)o��$����j��؊�B���Ҭ
�K�R��q�P��=��z&�2y�^��:��0B�<\�Ty:��qs�Ҥ����߮��qr����Ps�����D���`��mFD2��9�d�LLuh���)+~��M�(��A�Me_���n"�W��I6}'��k��TȘ!>Q{i��{!���*�f�?��9��
O�}j�=L�_43�r|iu-�sq|An��Cnυ�rڦS��3"*O�݋:��|��1���*��A_��W��#�`�G�*��Њxl��k�NH��A�����ql6��C�#�Wi�cy��8����N���f(
�Q���DT�ʢ+�4B�y��G�&m9���>�Aóf3����NڠMd\�- -闑��8Sk9:��+v8c�7���%w����I��VT�fg�yUM�e�C:�B<���o�#|Շ]�����ڬ�8�H�
�@!᫖�VSI^�~	)ln�>���?k}�~zc6����\�h�tz�z���?x�a�G�b��?Y;��k��*�2��^Nì���������kc'<��{pO��Q�h+}��of��KQ�����hz�?�u[�ܥ�	�:k���O�3�9&��5���@>k�d�����?;��[J@��|fU����+��CA�+d��f�J����A����SR?ɓ����7� ��̙�C�,Ǫ�[rJ�ʌ�������yK.��Q�Q\��O�$���K���q�O�wg'�����Y\��@^�M�?OQmA���"�B�;����`ny<c-�����%"��3�͝��`:������A�	����������H0���I�3�g��w��!�6�W�C�л�?Sg���-펬۹w���?|�C`���FȺԒ�n����mٶL���2]!&]0�g��O�t$����͡��Ò��������*�(@��u���IJ���Րj(�g��Mss��m[2��7k�ħ!ڙۅ�'�ϱ8�y�U[Y�wRO���Ln���v�q>�۱6l��k���f����m��j��Vm���Rq
�6=!� �5�F0b�cu��V��^4Tk~T���!���\$���?`�U3��e���߇�F)*��R�bB��yjL�(t@������㶮��i��ǜq �,��ſK$'��Qz�M =�&�ft%N���-W��3�X�o�o�u:?k��\A6��Q�B�a@jf*�H%��D��l�?��!f1�<� *rP��}<#r���ϝ�F���˰u~������&kzlFL2��w铣j�tp�cc��[?�< �v�>E�!�D������K���k��m��4E��%�̲��{�>�r���Y	���D��/�^�կ���J�d'���)5�$���I(��E�O�2�T�ɘ5B�`��F����+F�S!���4�o�8HO��ĵ��ѣ<�2��̋����3����5#3��s����7O=��JM�Hy�jү���2�ҥ��g0��Z?t��+ǲ61� g�RH9y��)�x�x�mU��a~:�/1N�qu�`ل�f��O����%���-����{EIH�����+#y+����Y����E�5��3���Jz�b��b6O�{ӟڤs��c�P�&�8Ҭ%�����<I',���؝�𦞄W�M�zԕ��jTc�>&�-B�p��T4X�cP��j6��Y}hZ�L�H������x�0p�E��C�Pe���cT�)������(�5�iUi���d;(��!��	�73�A�����H%��8��eDJ{v�S�	�����q
���:!:�jNQw&��!A���e����"�9ӡ�#������ԪQK\�#hGa=io?,$�Y���Y��.¬"�D��?���������V����.	�E��5����r��H��,������t��FR�o��5��P_rˢ���'#Bw��[P*֥C�`��]��!�G{���ܕH�4
ꑢ�j!�����R��}�s��嵈Q��2c?�;��$��'g�Za��i���_��kBD��}�G&XW�Hީ6���/�2�w�~�ۙ�$.
S���-/�-h�I?�l��+�j��a��`:/��Y��}6`��Q)B�iD!�|],ܒ�D���m�<L�AJ�آ�y�|+KÏ�C�w�2���[.]��4�jΔX��^�6�Ш�K\n�j�7\ޗ>yV*F���&?U�?o#:���[�g5]�0��He�2�xx�]�h��u�&Gf�xL���<�e�L�RÇ��-Df<Ħ��.x�LZR����Ƭ5��ڹRa�ȹlP��f��N_�ъ�dА:x��in�0���*9��Ku�B�l���Q)dE[�>3��MD��|G44�*
�gH��y��Ғ�8����?/.�XCG�yrG�;{�ŅA�=t�$�������|��_F��枔İҡ1��^{��7]�i�&"d�U�1K�l���(�����{����K\)�f�Nڧ���U�k����A�{b6��%ְ�g"�Z~B��	��}k�tbi���uG]w��ĳ�Ws@i ��>^��8��K���]Z��0>���Ǘ}Ј�����������P�J���a��و#a���2]��l!E����b�+�`v�ӻ��SI�|4k�&#o���J���p�ݸ�T�!��k�7ʲ,3�,򇢇31ԗ��!����t�� �����?��L�LC�C��$�Ц�V�t�$T��isGKA��)%�b"?͸�Q���B~�_
�A4>	�u�����!0���tث�zA�ҌCo�J?D���A�6L�u�Q�M^w�r�H)��j��ݢ��`�1�>��� M��
t��h�ۋT��u�36
�1�O�,|�O@K�\>.��E�m���<(����$�Ӵ�
2���"b�K�᷒m���,X���οn[>&���־#��>�bF*�k�\��+����v��J��e$�x�'�R����v��E�n�[����I!`&����Ko[��4Ϣ��O��8�E��C�3���g^hGd�����j�9z)����O�<�Β�n}5k8CZMfѤ�Ȁ��`��̣�SH
���:"���z�����#��RoI')�y�IB�fڙ��3LI��r��L�"K�n�B�����D�W�;C�RVn�Y���S�Q�U�'���[�o�z�ޡ1AO��?���$��B���n�8�,��J)X��5ѣd��wݣ�Jt��V�zJO�����u�|F�P磞��>��}m�p���?78��/z�9�I��N`�H�'����W_�L��.#�\x�����ѭ�Ԏ�T_��o�m���;��Z�ja��TP��x�
�h��B[�	}�*H.��gO��n��9&��E`Ʌ�*���Cʲ�>�C�rM�W��2��O"�����[@!����T�Zf{��.s�,�xz�N)a��Df(?��7^�sF��G����8۩�g��c�<aw�h�e���ݮ`U����2���[��H.��/�&���]��f:�<�7� #����������0իxF�Q�x�:U ב&;S�\LӘz���.L�xWW	����t�dW�?2F��\O%˕�QpV��<�`�6��+��Eq�������
��X7�co�C4�^��J��7nİ�3���2�'�Q��ˣ(�ʙBÃ�|�7A��A�ĝ>�|�LWi����.�<�9+/ *�"\"p�/��s�y-����s�T���x� UX�exS��>l���K$g�^��gH��%i�⥄�<��wA5�	�n����x(>
t��J�4�H?����T(E]�84eR��;��`b_�}��5?��$�?e`����8��HJ�9(�6S5�'KQ`��	�2����F'^�x�G���J�D�'N҉��3z��o=%�d�>3ck\>�wbc�Do�Rs��sQ����[oP���lmXP�u�C%�L�򼘙S?�.�!£�_G��Q?�� �V�x�@N;Y���%a;��H2:�=mHt �z��	�UU2nH�0���D"�w�,�����tX��Z�̀�cثޭ����ߩ+���a99�_�n���g�9+��1�5V��.�p/����| ԒƮ��|j��b�G�{,>*�#p:g�a*x��d!���q�?����B��ΐ�0�Ԋ݇.I�'Y�{$�׆��j�~V���\��l�%B��8T҈�]��~�J-*¼�a��:x`�x��x��b�v	�^��e��x�+q�K���j0J����I��V���@[��o�[�������A��u�v��^�]��<���3�ӪKI�S�]�z��3IǇ�Y� ���>�#B��/9����@�.�Y��v��uK�y\q��?����[��<kpu��`��ۏz�}�eHE��H��bJ֙�m�Y�)Q�I�tב?��E|�bB��.�J�9&�1��	��QӤ^��YCur�@�D�Rq�K��bU�WJ�ϭ��Of.=�EB;�kK�޴	�dD
2���e�~2�ΰ�r_ڡ�0-���p�>\q�iZxO�N�.�Z��AqO|����'�C|��rf����a�J�DG�M�0�TR/lb�=[oBTzt���U5 k�
��p��1� ��Gت!N��ė��=q8�^T�Q�B�OX�vu�z�ߋS��mp�P���U����jJ�$����w�����]>=S?Խ�}�����S�RЂ�ވ@%rV�����t�i���4��hQ�݀3��\%1u%j,����ց {m���jUSL5;���~�jJ/\|,��%��z�j8ܩ&��[�n_��[L_�D�@6PvWC5��rc���#�h����	S�p�$0,�`�e~�5-�Cm�nG`��V�ԈEx���p�������R���(��2�n����7T�p�+���F�[��䔋J���[����o���x�Ҥ�rl\�S���������æCK���Ѻ�k4�F��'�e�ah��A�QԪF�Ư�Y��g,<na��g�f|57B���k�4uL�lz�Ɵ���{�>ۢ��sq�>�c?3�B��?۷��Ǭ3�Q���;N��	ђ��-��+ OK�/��w����11m�ֆf�uu��m�4�<��J־�E��x~�*�j���w�u���#`OX*P��Fs^��NK����{7�*)#�����'��`� ��|U�JA��"u>R&��I֎e��Ѕ:D��9/�D�b:�TZ�R�Ex���a7����E��NsH�}z�R�+X�"5]��=�t��`���ߖV	 �!ǯ���5�0���8By��Lਇ*�~$���&$�Ҏ:z�P��~�����|��\��Ǔ�*�p4Vr2\罹v���g`�􏯎7:($��p{2�k��|/!o|��>Wۃ���5}Op�|�//P��0�tɃ�6�\(��W�ݙ�f1�()����xZ�4gT���Ћ[Ur��S�<���� �_��Rq�RԔRTPzʍ:mC��I���v)yt�h���r��N3�[�šn
�7�bS��UPx��R����<�ƙ�>�~[4҂��\	���I8�_z�T�z'|o+�[����)L�=�Y���Lꄽֈ�<4�Q23:&�=�r}]�}ؼ�@m ���x�t�d���g�>�J$����ŭY��C�R*�N�g����T�#}��ҍ�?�"^[
5R�y9\�����������E���(���A[�vj��i��[���h�nv$��[�x+�������7�Yʞ�bW�EK]�g��梽0\�`5�!����!�'�b�������,�y��gĭ�KgMwۿՏn׈>��8'�z��~��4�|�Ц�_�_��u��(M��ЫUې]ʆ��w�9N�m�p���d^xN��8v-�G�oχ�m����9��^*�֋�/)#2g�ئs�a�AU?i�-\�N��L��$��š�c]�\�n��b6~;�!�r���F�����eCZ��^�
���6fA4z�2�w����ٰ��P.L���(��?�D�{c�o�C�����(����x
���Zt��P�ה󨮺��Q*���x�����X,�TlӃ0���Ëw�%
��V��Ǳ ��g#`���'g7���#����$C�;qwtceտ%.y���o��5��h�}%�6ɭ���~&�'���j��V&\{$�)&�S8-�M���U�G��O51#��Sp�~�?����ߢ�fڴ>.�6&?A:�x$
{Z�"�0�RX�5��q3%��Xθ��Wt���W��`��s3Ka��d��
F��J�0}�5������+G���� ���!w6���cݣ���l�4L-j�n��vF�Lu	����Q��N'���-�}c6�[d�Y*����.��p���əp��a����8m׽ӧ���1�a�d����d�7�夷-����Ѱu3?�����ɢ��%���L?U�^�#�D���F�aR�[=�y��d����EbL��L?f�<�k�!g.�����I��0'��������xT�a�/�_������ϻ/�E�]k��]�3p7��3�JS}��7���C�-��.+��9�$�mX��.���7A��)�F�?|�	G��v��-���/SD{-Ŋ��d����#���.��D�����`�@3���6|���P�y��闀k�Ӑ��:�䓱f���]���g�@7>q��a~�f�m*F ¬���~*�j�ڠ���q�^#��C"�m���*���w�ڀ,<񀷰h/D�ʗ}�N�3i&�P��C�V��A�L=W1���9��pȆs��}k����u��y���g���׸��*�6/P�m�>��<�#]����5��M����=�L�F%�_S��%�֚xM|���ȅhe�R�$F��G�Ô~zXX9�|u�b���#D��-�w��/���u�QgْՇ&���w�)���Aو�ӊ��a������X��������?'�»	�r�=�
�$2�D�s�s��P�������P��)�g��-1�A�j�v(��+Q�;.Q��"l]�
���� ���5�ޣ�aF)����@�]	���&:��Q�K#1�����!@���(i!��>ߞ��n�K�Fum�Y����[j�u,aӈ���9$T��S鄮��]~x����B�C4&���.Xu�o�p'E�� �_u�yG4��]�%UZ�Oѵ�u/���(�ε�ꏉ�@�]��
dL����δ�kO%C�m�~K�z���/���Tv���-�2|�cvk�p�t,%٦�-�0�oԥv�:��ӎS����*�AY���k\��8aJ`�ZA�2�t�2(
��4L��p�ͤP�Qd���~c2=I�G�	E�P�1� ��F���Q��{�9���D��`F6Mj�@*��/Vr��7׽�b^�jH�ȪP'�@(U�a���4�>��^�]��#�N����gi=��/��͟�+�-�KU��V�~�4�zcӎ6��\�S�$����7�Y����bu��I������J���:�g���f���D�&8�.� ���=�����J�	�q֜`!|7P��{+=�(���-������r�S%�3l/��Y��2�o�@ts�ӡ�p�^�*���`7��૑��5Jl�(d=���$�0�'����	�@B��r?9WX噎���;+��&���V��p�� 9�T�R>,oP~O���Q=w���(�_�QYBAY+�8�-Ӱ=!�R?��I"�{���(��t��ߕt�]ޡX�C�#z�,����<K��<N�M&w	7�؃���O���B���9�	χ��Rw�"g93�g���s'|IN�F�Ű�� ���}KM�"���N�������߅����_t+.���p.,͝4��t�)ƍ>��q�$�����fn�{�.{�]!z�\�>-�UP�t�r?�Y�$殸f��ޡ�g\3�C&�m`�yV��H+NS<�v#�LRC�M�Rτo93�d�/�;��E�d����7���#B�{Q�c@�%�<��!ƺ<�ڳ�}�C��y;�(� ��6X�?�?&�9:��6�ضm۶m�۶m;;�ضmk��%�ﭷ�_}�꾧���U��n����,���qH�L�[�D�3���k�H��!.�Ȓ�� �onـQ����%eoj��߉9�d�:�qi㚤g�G=��+�c�T���c�a�+u��n����[W��~j�Ҥ��/�ܦZz���n5�i9���j�L��r���2�u(�Fr]�/�W$l�������(O��<�}Aq����D�����=b]�nPE��qit汅F�����X����l�z��N|g��٬�Ž=5)?h�~���۪���?��|�Ҙ���$F�]������F�t{"�C!�o�*D�~�>H3�y-� ;r����~,1GӅoC�b��:+��ߪhF��IG�1��20y�,/B�T�qQ��ZEK�it��ޒܼ�[�H����������������	��1y���''�M(�����S��,��F�e�����A����ůȔcT|Q��Ԍ�
we$�q�1��f��� i�=���~�C��=��8�U�6�UR �`�l�o�`��gN:gR)�q&�f�3�t�y�����\t���Zf�=.�|�'��� �дB��t֬�+�P�(��᚛9~���'�����h����{�����k%<��Z����e�k�cv>fGfTs���V(�ꕢM�n�@�P�*�y��w�3��i��C��;��u>�<d��羞�$nw#�tw��@\��Kow���m��U�`��ރHJ�k`T=a>����65]��O��c�+y0� G�0FR�����ޥ����S�Ɏ>�������j����9xΗ?�k	(��o��7���c�u�o7�g0)*^�T�X���篓Q]�ڡ�����(	��2�����"��T��@];�Y�*ូF2\����-��.�2 '˂�J�}m��R�����VĶ���D�'*��~/0��;��=�VpĎ�/�BY�������}���k�sl�6�B�h����Zn�KSLA:�N@1Xn��-=�zJ��Wjza���]̗�k��D��ـ�!���[��CH����7��Q8#75�K��a_n�-T�:sf8K,ٻ���V�O\�@3�,���ﾴ�Y8zv�Q���M9T���p�B�B��D�&�;��\�oޛ���/I6����d�}�݈d�i� Z%7�6�8���=pviϗ��Ui�OV�{>�͝Jo��k"�؟��/Oݗ�#c�;kY9gKy##�����L���" ,���+��SGr��ۥ!��"d&�!��핀��q��#B�ގ`���.�����~��]&B},oy,6v��>���5/W��#CG��H1D��jՔ��ws�dG��2�I'%IU�l�K��$��XO�oV˔!&j$��.����:�� <M"8S�"�1n��C� ��ʘIqL���z1�\o���ky�a�8��k;Ux�.t��Ҡy�4q�.�I�+1+_�b���=��ڨ4@�h���&#�B%^����w]�=������M�y��6E��tm<��abEo��D��3$�0�h��N�B�d?��sܘ�M�����r�'�L�c�Di��JI�sQ��|bI^ឦk[�4�!v��	{����)��Q:�feg�j�X�v�D���Hqv$�M��ޫ�v8θ����`���Ŷ�A�Yԃe���e�n�E߈�r���Pft�
�#d�yj% g6���Z2(LQ9��`�����Y�q�/�9�-���1@��&��9��;�5%��~�Dπ2���?is)�� ��q����]�pZ�v�w~'0�H��Z%�q�����)��xH��I5���Ƕ�2m��V�zZܹ(h�U�ڥ��8VX@$�Ѽ룦���b!�1:+5m���;v�H6?��k>9�BC��	}�p�al��I���h-I7���:��N>Ҟ0�j�\Ӊt���g�Ѐa4�$����|��]:Q��Nadc����.�)�nj-��M�W���@��L�0�[NZ����0�q9AIЏ�n����I������rՊCH=�����X�}��b!�mş�0�AM�U�������1+��ɥZ��ʼc�&�hR(hІ*C��"�iG����
p��t�,8ʄ��3�P���_�K�-��"��~��W�������SN��g���N�s�gfyY����m��Q=�����[E
e&�q
c��q���������E��|���j��+�A���������N8OiV4� q�8�T.ռ��C?\7�9����nq�[��@����b�W,j�'��eɨ���[s�š�'ѓ3s�0*^o�Cܾ�ѿ3V�Q��'M��X���t�+�(�:��gy�K�>kAu��4)��Z��J=E���t��������%�O@<Lq@�'�#������'đ3B�XC6\T��e^m�,��� 'Jm��*�N�5�Y�b
R��_Ƚ�F퐦5eTL�RN�0��dku��<%��;�m�#�.1�P����4cT����Fqz� #�6*Y�*��P�kq�`�dTC~���.#,�(C"�8���ך�K�����ݓq�'t�{Pw�_��7ǝ���b6!�G��J ��8U�R>�*�YG�1xFQ�ZYY�Z��S�E�U2�˘	/AL�=n4���#p��H��.̛�Ƶ�=~­ͨl;�e�%�-(
Y���[�X��c y:5$f�B�dbN��(7�u9R�����p�5攷�"N�

 �*{Z��qվa�1��*&mu7����Ph�݀[�`��{:�����,�����B��Y��Ԗ���xu�z��ܼ��!��^ ��T��(�('��gM� O��S��a���il�x.T�r����Y�����Di�g��e5�|�
�d�f�Q9`1�5*B F6ڏ6!���X�4��ǳ���h|2D5r�-0u��[��]����G���`�=�](%\�רު���$N
�����*��G�4K��K>��Q�1MW(b��""O�#��HR�u,� �Z}�~{���|_�¨S��"��u,:��*�r\��S�����ĺ\~�e��|�f�˖�<��	���e�R��m_� "�EC� L9��!m`�*�Ǧ���f)�]�	�[!����V����}]�s;?D�'L�H���Eɺ`'ߓ�/�+s6(����sLC�&���\���7�EW�A%(���_]���]t/jN����kty�9���������G�F����u1��xuDڷ ��W�A8�<���'q�-�Β�V=�L�q*�`T�10`��g"1�c?��r����Ո�\�Pk%�v��dh� �	�V���-%BG�t���N��������($� ��z�қ���o������0J��S{ߢ�����c���~����a�V'�I�׹9ܝ�ð�����_�Q�g�rɝ�+&e����|�F�)`�~{�V�1"+|:��gu|�m����r��v+�u���.G�,$`�F�k��A�jE3�{�,8h�C��XX91��9?�����B������s�G�^Xem��J#�r��n]��ψ[r7�WD�{����@��sr�ڲM2<��t�v ~�&،c4g�D��2hl�Dn��Λ)�I,C<UC�,�����PĔ{�[������ ��宷�y�<9is6��5�j���!#z.�M<V*��������C�s�F+H��XD�I�H���#L�a��<25,��6��ṫ�>��ϊ5S��X�ȵHk���o1�ySO��6h�%��s���D��T(���.{n�v�i���{�����o1�Mt���A��KN����xM������``�N��gW�dا���Aϖ�h�ϗN�����)'RZ>:8��I%�d�`�Hm7���xI�x	��@��1ǆ(�c�� �PI9凣�d������Rh��#�m��M�_����7��x��Ls�*�𑃊κ𯮣��9�Q;w�	�����tF�O�|��W&��5δ�>�H�.�rBHL�/��#.��,�rH�*�j��~��k=�~[��3����b�sn��$� ����q��p��%�E���=��S0��[&���?��S��K�C���!�+��x���ղ\����
#��B�]����(	rC����gN{�R&�*/Sf�=����(�oG��-F�VC���-���7ש��6�"���z�~v�� ���g���Wv�����:}K�e��M4��������R�:�������(���Hi���GR�]Ѿ�ES���o�F���5-�̟Yoq�j�ɿJ�ԕ���/��&7ת��;����� ���B��|��ܞ�����z��^����e��^<g���� ڴ�����U9$h�@��G���ӏr�ODEy�3-��O{��[����I����rۥ#�U����+��-���+ؿ�/EP�vG�<�`&�#QD����d��Hf���4*�	r�h$�`�ic	C :V���iz�K{���nk8޿���.+�c<�=M� �?`�2"��{���h�穵�����Vk��G��?��ė�C�¼�M��!�ܸAJ���ZˍF����3"_��#�+$��KG��cfx�+R䝏&�}�vX�cj�S��4u��~�.�O�������!u���S{/��-7�����S������F�̜����	PsG{���P��K��2m*?�_�<p#N�'D c��&u-�;26	R>ye�>4P��3G��S%iX�txz��7����&��.CX���6��5��
F*��>�r;lvev�3Cm��@���@A�X�x���[!}�-����+��S;�IP�S�,��^�vv39�o�pR��3��ٲ��DX�VYT�⋯tB�������\9f?�>#YЫ2HXӚƬ�J�[86����Q�>��A�k[g���l�,槂��(��}��\���=L(��Zڇ�z��~>�^���v���`��p��Y���	�@���)����S�Ad�{�\�Xf�
mj;�||�����&W�{�g}Sa�V[�6��*�r��ըz�֩JbQ�I: �X�1�v��s��{9�����K؋�	f<�C�:&�z�tz�6Dl�2d��b��,`X�ܧދ�~��у)Y^��t%���6It��2? ��lP߶��ʛ��	���_��~"7hh]S���(��ww�]�{a@�� ����C��a�)aŰ�j��;12f �V��t_�d���s���CK�����U&d2��y^�w��îȜ���ˌqQ�p!�)��U�%�#���G֬|��&cbzy�@�1v[��d��,�!�������4��Z.ױ����%�H~ �Ԭ3�Xc�^�N�D�=��_ë'�P�֪�4߫�� h��I>��a�#�N"Ƽh�t�����'}��UÆ�s���̕g��]�5�i�*O���0��>0��F�#�`��\����/6�)2(|��{u�_�8����}���~ m���#����BG��x�6�~����K?���q�-h�4�g��WY�f\���蠗K�r���K�vt�)���SR6c��ӛ\E�z�q]'�ŒJ|N<�3w�}kƼ�'7#r���Z�s��3�S�b�S׎��c�k5���,�
����m��^L=\���K�(Bi�q��&n/{ˣ/��)����#Nȕ3���^6 ��^2-��.�ר�h$i���~��D�~�:��'���a@y�u_�C1�%�`#�ɸ"��#/MjN��`(�I����9Ҋv�(X�)����o��銃��i��#`|��ĺ������D ��m�*�bR�:����>�s㥑7b�\�CJP���9�u�%�^��Ѵ�G�kԡ��jD���}��g�. �\w�I[�Ҕ���vS��`&����4�~R��W!���r���DI���f�z�� $
�ǘ���P���ϵ�?��s���b����I��-֙�Yv��9�
g��H��Ŏj�sA(5'�'�Ux�P{�-�V�j/�ʚ�ƙB@gi�<���}`n*K� im����S�4x�!�n"��wۣs�5ܣ�ܞ��M��<�G�[���)n��9:F:2��k�h�\��ɶ?��-�Ƅ�сL����|�2N+Ѡ��KI�����:���㭪���co۲�me����@]Z�0DYOX5���
���NNʰ�$�IX��8."qPVn;E�OCQ��H��p�u�)L�1�NicvU�����7+�5�9��Q<�#FM%$ƖJ5�3�vy�Ԭ�ؗйPy��?\�3���X�<E6�k��|)�ى��}ݕ��YA��p觴��R	�j�����9����C�;F�i��
l�<x�:�l<_ˣd��mO6��N|�����F��w�Ƶ��'�/u�(���Ո�ۮ^�[��@G���o$�I��<�RX���z<>ʤ��X�}P�uC;��t��d!��V3���e��Vj�y��̮yw�8�?����#������ny�gg�{��I�1O^�d�u�xx��<�<��2��5Z���� ���D7�� &&�r�S������������G<I|�z��)5�l-6so�+e��4T0[��ġ�ewo���0���*_���Ӥ- �u O��8���Xr�ꏘ^���Z�f_�z������V0�P�tz6o�P���0�2r�sˁ\LR@9FY���Y~�p�h�Tw�E���h�#�I�D��rd
�#zpz��UY��E ���Ю#稖�6g9"?�cQ#���a�F��l������6�N�i!������I��6�HD���+,5/��s1��`�5�@��X%�3OaZ�a�9�S�[T��(�4O[{AOr�3�U�v��q�N�#%"j�\1qFRH�����l_�ֺ�iUə<�{��3=!~/%�=�zl��ꪋ��A��������o����_�����E�ш��B���O~��N录�ե2�u�PA�Hc�)Y�'�da_c+ً�Di�]RsG����b���n�G��fV�#�m}�	��t>$a/v�69�X��#4��#�SRC!�,��_5�6=n���Z��"a,�a(my7�y���㲵ۼj%@ķ���9L)�����_�����L^��I��2�úe`|��%WΔ���tǞ�P&,�p�h!%aү���nq�K�Y�w����E~�M�q�H�,�\Fl�/���U\d��a�����ƘҐ����+fb��t��Z�'^� d�> b��p�tg���69�,L�_oA�O�0���,��,,�w���Н��A�fᶹ��:�-9����N�� Δwp��m�Y�>�dIr��)�|JE���Ysh����s ��b1UKʔ��D�9B8���wKry����O�
s�0�]����*H)qLa�w(R�n��6� -�f̼�H�,��W���v�a�m�Ћ=��tJ��=�1�5r��m���� "�2����Rz�H�g���ZJR�h���`�J���)���"QS� ���ׁ(�l�E��H��_o��[w���4�b(	�'�����i6�;:*�TAX+���Ȉ�&�ɟ���\=��U��x`\�x.ȊS��BсR�sT�f���������WtT��N9*�v��+�j�}v;Bq�nIA_���v:9~K�����@�F�Z1ĳ�
��AjH���|�NT�t	���w^Ů��Ns�rh��JT�ܧ<hczn\���K��A�_g�G��KT� �[>ET |���YV�%�&�A��hx�in�e�͎�@}�F��[Mo����o�.ޝ#h�t $/���;�F���w"��n- O$K�^Zk��_���Ӣ�C��k�@-O�ӌm��K��P�-�k�+)�.��_��B��`�+���it�E�P���pP�{��L���Z��E�Զ���8�
��Ц���Ǔ�T�؍�A��owoW�T���R��(��N�l|;;0j/�8��d�Yw]��#����u���]
��$�~3V��ڥ�|\j8h!��F�G�/=�����M/( �x��/&�k 5=^�79W��"	:�B��<<uR�C�C���&��#$�'��b�vo�J�����m�B���߸�ё$E��)R|

h�k�GE���8��z�8��#�*��$��e^3v�|ӽ����m_/�^GK%>����J��$����E�vW������TG� Ģ��IP��O�A�]f�M�s�ûrN��w�1�Y��J����a��t��]�ݨuM]\�DF�x>�!>�g+�%����ʬP��ʋd�{�����.��Ft���W%�0�,�i���2&�E��Ƒ�6�VL�O ��|AWL�Q��8FH��� 9��\�B����ouMP\<��>��r���kfbe�M�
�[��%�MK�UU���^/������!��r�D�k�M�N��{n*�El�B�
bgD�V3DT��LJ�dt8l�-�6ۗ�c����].ԅ+��e�����]�l;�<�)gͳ�Z$�7g��]�7�j����g� 5�&��
�����zj2c�MX���osŒ���0�H1����`�C��f�Cn�%GC�蟑N����aX�F� ]�J�e�c��Ki� �WgQ����]i@�S�$�A�9�  ��b$N�������ֈJ�0/f�����UϺ50�i�r6��ީq����iV�=��'�	��]��]��;-z���������a_�n[O�o�I�{Q��Wۤ�9o����\Rufc�˦��e�෼]�ؑܐ��$�F�f�x�r��'�=�M�s��9_�6(z�܄��v��;7��넜g8l)��%jc���6��c27�կ41H�-���%�_Z3���=4���4���+K�~����c/����@W��^��x&L�)�a[J.p�b�fZ�-�C�?�9�*Ž�Ff���f�{���Hnż?�T{���Jo�����1���v�����Er<Α��<"Oh{G��Ub|8J�Ʋ�5#~�I���ࠤF`K8�g3`��w1�-
!��˶HMhmҒ]�D>(�`�p�q�K���������_�O/���Y�o׺��Q�,V<���CY�:�CB��B~ڜB��'`�幤���._�8�a3�	����j3_�0�&�r�u�ph�o#/ؤ՗fX�%����7�y5��S�`�W� (�3�YE��J�l0H�K�f��{ pDn�T�q���_U����-�:3+F���慽�p8�5.o Qr��9䏰*�/F��| �i9�A�J\l�f��x�MU�7Q#Ƅ�K�P}���cmA�^6��X!=5�~�#l&�\M
p���}�B�lJ�{L�/��H�Ƶc;SUf�,ޤM�ê�dW�r�2D7���ۓ��C���Y��{{�x?g@�0��в�!�� ���ۃ��l���Y�d� �ं~� �@���"0걸s��ɨ��ٽ�Wh�$�8��G�L�)�I+�2�_���w���i���ѿ���� �=�W�0CeR~!H�lFT�쩱'��Zt+i	��D(-5�*��K�~�16l/���N�Ha+�$�𚽳4�"a�<,���2j���P�Y��j�!1�0��d�q��4��kЅ��{��3'�Z��4�����,<�`��G��bU ���О*l棑>I�f�s/�]��ʤ�A)�W�0c�L'X�eЪ�US=<�ɾ+�G�ar=`O~���X���H�X3!U_�$����2RF\d?z�$����L�O�@³��d6�=u������C]]���o�������լ~$�.��"�����UF��&��\�=��p��U�n����{���Ex$l�P��7$4��p�n�_:M��T��R\���۬M�3FT�n�}��)����O�:����<��x�R}�[YS�o����ǟN�%����,�$;��e�� %�&[-��k��`%�K�wg��1�l<�,��Z�
��x�Ur�
YHEr������#Ւ�ڢ����Ł�J~���p���x� ,L�R�������~K�xH����!7��(�7"������`P�� ��ls�������X�9R��k��T,�U�a��-�X~!�%��Ѷp�4�~�=�.�����2���ARb�QS�ryq��\�2l\�3��Թ�B3k.���t��iB'�MJ��#��{�Oc C���(7�a����~Hp� �8���q�W��gi��Rۜ�Hڰ��Kƀ�Zt%����oU�4�\]:����H&u;�g�w��f��������Æ~ğ�k�R�0�,���_RU^A�#J��~g��5�$������-N^�/w��E��_� �T�?$M�YrYī�@��#���]��,l�Ce�~��- �f"��DA	",?:�@4o%����"]۰3��b���B���f���P@�/6��9-y���ц@�C���Fe�����D%&$��"ٖ�-^^���.�X06�i�(g{�>upNy���;%He(~Ch�������G\�����S0���,v�LnNw�vbN�k�C{�8�l�Q$M��G��M˦��z�>�
���o:y$=!>��6c�y��t`=T����x���7����TZ[��ےZ���R�!P~�%S�E4��*r:b��?�-w�w�h���挠��Xr�L�Ɉy?p�:��&D�(�4��;m����kW��	�a�
��@B�5r	��NK=�g�-����w]%j^1�0�W;r�u�.X����#���˔���?�:�x�g=����Y�v�3}֞�0����N�ܸ��N������,�6�c�a<(b �BYbB�7{�q��~�7����MdP7nB[n^�Z��in#j�E"���A ����>l߽�u�s��0��A��l7����M���C/e��}��m���VP?c�V���se޾Oz}d�~�m��s���W�w�a��È������`�Ȭ0o������3���IQ���0F�"� 9/����p�+0��{��H��V�A�&��\��?K4�p�]�;ٽ����'�u�/�!�mD�7�D�W����y�߾R���w�X�~?�{���b@e���������}���j�wR}j�U�边��e�l����07k"����C����Wwf�F ��9�1��g��g�da�qa8�5[���e��iF6�;cM���n$u���^�VI;˜�,�*f�~1����M4���qN���bdi=�꒿~*<�V����\��˩�Q$o�X�X)
�BѾoż�P:��?"�2���`���0����G$~X8��e4pZ\U��9Xl�}U����G,�Ͱ���%�'��7����ťh�$!<�&�2�Nx�b��q7���2g*FB�
���8�e.ܙ���������^�^�(f�`�SW���v~΅��T�9���΋]6~���4f��}(Xլ��o���<�3t3դ��h�;����&O�ⴍ�.�����z,��T�8�8 �<
(C�g��'NK(B����M�OtAb�@H@�'x�ϱ�170J� ������Ju�6P����н,�Cq�����G���cZ���E����u�7��b�J��x8�T������c��%�&l�l��2��1��Hə����v#Zx���&Ҧ�W!�P��(����;9�Kˠa"	��ՌD9@#��h��ҳGZ@��.!��'�H�5Y��n�3+3��A���6԰���e@kjR��A�S���w���
�8�2ª�ϸ��<'���[�o�Z$�ŽMB�?f�@�t�W�i$�7��s��9�x?�3
ʙ�+�]�m��=��ͅGUvi��67�)bz�%nG^�@Bπ��^Ɵ� �h\�Dz�c-��v���D�

�ɥ!l���/��vÜ7%[�6���G����k��/f�ǂ��k��*��悲�~m�ر�g�3��*���H��+j�t{�)��v�Xgxf����=Z���,�
��H`ξ[���nv3D�e���1��B�\=v�����V
˖�?��H-q���,fg�	�ф]lٯ.Q�E�+�� @,t޽M�,��xH���Փ��|�`�b�g �an��z�|H�S0�3�/g�nW�4R�!�ͺ�ɢe+��@�덪B���{�6gټ6ohj�kf{ߥa^��/��C�r'(�$t&#���(K*���qk�y3��t(�_t^j6m�8�uj������h��2	C\%��A�"��� eŐ(w�����K̅�ˢg
g����6���N�4��>�����y	��V!���.c��^AJ�_��q?��
��Vzϋdo"7�w��+s�/��캛~��ӑ猆�77��^Ϋ�iN�o�ߕp�eZ'��S�:���u0pċ(A�s�Q��b�k���fD�����T�(42��eT"2�����ұ�;ۊ����RNp�y`��D/��Ɂ�kP��,� �J�i	���r���g���a�r�5i7�h��Kk��iK��^���i6���K�nx��f��Z�@�̣ɵ��i�f����R�Ķ_n麗�Mn��U/�x��������ە������
S�b�8�I�٨��O5�Gp�pF-^f`���)����ezP�S@���EW_��9�q����n�u@+�2�p �����`(���|7Dw@<
�`�b���z;�M�h�6�Te�z�v�4]-�����5�
dN�=g���<C2)i6yҲ�$�7�m�,
A�d�%�0�e�9=��qs�0@FS�O8z�쮍��#�]�A\�MX>��%7����?�:}n�Ɋ��б#�T7p��vv�
!�l{�����F��ȣ]>�3���J�E�-��^)�&7Œ���J�w�4���$�g��!9y�@�f��e��o��M8�d�	�s�1'�j��$"7�M�l�Ē��M�-{"S��MO ������T
z;���j���J"���z>,�`_�q��%Ǥ��I(�R���{�֖(\Ǆw���M�����Ͳe\���H$ �����u�l0\�)����[�5���hUP,^��Cеm"�Rp%�*?�d��<m�U��\��؝�]�C~ZH��8E
�UsEYqy �5���Ib8�]nh��i�مð��vE�K�(��`�����z��y��?}��i�51"������j^4s䔔����gU��V���7�zB\����� %&%;�,Z��
�IQ�QR�^���̲x>)���cx/kZ�^�߄�u��=�����~kBi���[��XH76\oi����Z���s�Τ�P
^�<ct��+�R�
���F6���4I )�C�,���v��arcI���[��/�n`3O�=�hs�O���
�[O��/Z���a9�Z��1S;I��s�^���r��fY�$9k^��	��D�]��F}gy��01׬�_����4��?X�JmBU<�+r�>�IR�S���K�p��덣X��gn���i��5��8�XO?]{ܸsjܭJ�zZ�8*�g���s��Q���wjX
���JZA�,dC֔��ˆ�NPQ�Dl�J ���]xpR!=���.?m�@��,��L��]����B���-L��1��q�O ��G%W�P�^w��֟?Z��ïS�L��
T�����e�l�/�V�*I	��ϬXE4v���Ꝁ�U
�A��ڔJW?�#�UT-JR�(S�`k8����y�YvhE�Q��J���⡷��+�������\V׆�_+�"K �R�ݜ�5?�T>Z��Κi?}z���k���+��;��'���;�3�C��t,���0"Vg��W��2ϭ���u�u�����SRQ��d�u�#E�|����GΛG�	ܟwÄz�밑���xm�{�ޭ���������(.�Z���ئ&J�'��0_;Ĩn�Qy���X�]�,�Y/�*�>��xǧ�LD��L�@�v�^�&4���K^��%b!�:�|��f=3��7�_c#��$t�����d�4�.B!)���J����	��i.�/'As��q�)�V����Rw���tG�E �_?5?�f5g�?��n��!�?��^���VOw�W�T[cW�!E���z}��x��J��z�LS���T�s o�$j��!�ܤ1zE,��q�0?����4���k�<��25zy���޸��ۂ����h�!u���T�/BCpD׆f��_��-�bE�fO�<��ͥ�
�p�bd�F!�����T̹���E(~�h��Vx�R�k��޺l��D��C�6��5�	'���Ͳ67ͥ���s�L�M5W���-H1��qo�m������Uo�I�u9e������9��AN�:���&^�Kk{���G�����.Q�dk��ls���7�Nk�9s��dx��N����)��xpޘ��s(�� �����e+��ۚ����h���u3�ܕ��_|��J8*�/��<���=94�ݽT^r�������sy��"ʲg�H���Q|o"IJwV��K�k˪$g=�B�?-4�ɦtx�C�;�om�>���[����uQ&�W<Tuӗ}/x�P��,�G���˺/�*����7������}w����Y��bGrW���ˬo�Z����e�}�_=���r�_�_��'8���+��
%+�����lev���=?��=}�r�Q��QHc�,G���iħ��i*+JҖ�t��Br4���䋴{�\�a��~6��5hyӻ�O��B�.LB�� ����s�3 ���uIS�����*�a�B��W�1�Jk�98��ns�|o5�<}S��*����ͩ$���ߵo����EF���[�fsX�&�"�9򔗜��ⶀ��Z��C�=�/�ۣ�4����Xk�߫�<���DT��)�S8��I��i]7.������>)̥�F�
�fJ� �����/(�N��ߙ�@�S�7|8�׀�F�k��t�Gbj�ԧ^g��MAw�\��aԦ��d�;��Jz�̡�?�nv�M_ ƞcE�@�P��n�E���R.���m�S(�ʦ��/���~�����ER�;7H66�o9e��E'����(��k�M�@	���:+���Tvyt���n��N�o��e6��s6p"��	�������g貼M[B?�+\�a)����9G[��e�0�A.�y��-�q2	�W���x�2P<ݭd�m���ɨLv<3٫;O���E�&ɹǕ��>Їܬ)���鍣8>��L#y�U��ǉA��܄�*�,J����� ꉱ�w���?�vw�=u��)b�;ܽ:^.h�dUN�/��g��~?pY ���b��s3k�e޹��8;9�%���|�h�e�AG��]ݮ7���)�ڡ�Q�l�����扴~���wF��K��Փ:ImA<���w	��&��{`_^~�!�d��DB���g>J���Hqx}��h�5m�i����:�Ξd=�J.����	CX�^n��(=�&|Dx>�V�oYY��ߔo4�f��S禁�3�R�1��k��f��܄���U���dr��0��zb�a�o�R'�4A�����Tc��.t���^$�d����s�Y����r#���]*M4�b��E; N����0P:�短����y�4EƆux�bF�f��@��6���rW`M��g�%|��N{����Ō��#p)r�o"-P-�d�~{M!���᷆�����u���[Qd������sD���ԸwE��#�?���HZz��e�����#h� D�i��������%:�8ߟ�n��dD
)w�+.8=^',�UY]�M/�D� �X	�߬qt�H����ld���˻UX33=��v��oó�~`��
������ʊ�����ﺳE�QT�G\����"�ﺏے��멧a���'���(��O)2a��ѥ�&����u��oG	���	/8z��H�f/^D8rJ�,�CtO6qݎ=��8pj?�e�]8��~d^�Mh���c�T&ٛ�Yz��NZ�h�Z��Ԑ���`��{� ����Z庥K���a������e��x'�t�f�:��w�ůH�_�Tn����E���.��$1�������8uӕ��7�����\6�����!�Ns��=�7t�Z���jR����QҮ_0㋄�8̲���c+��ʋ_�5�9��� *H領��?eF@����8=�PT�z��s�O�QC�D�`UKu�obJ)Q�W�p���0	����]A���Si��u�oy�X���[�.q�&�+e?�E;����a�zBI2��T%Qh6z�F���do�ƃ�@!����V���W���M��*�>/���=-���s���i�ủmN�m�Ll۶m{b�۶m;9������������t?���F�ӛ�>�M^j+��H�dX�*��D����P+$$*��ힳP�٧l@aӭ�%M�yBh?�,w���H�Ԣ�:h��|�Omr(��-s��Cԩa	b|�8�����e��y�D���������0�V��|[1y���Lާ���Ck����I!�f�[�ع`#׽B�KL�UB,�H��y��(�C����Z��p3v�ͅ�bIr��_������Gjp��>@����G��f�Q ��	�m��%�6����?H�v3�����ϷV�M|w`�Nmx�iL�d�!~H�s�8?0¯��ĥ�O-?ǲ1���{����*ݱ���Ert6x}�p/[��V���X���[m�jX�w#jӚ������N�{MZ�:���
��mϥ�G��~r^.��/E{մ����Wɋ��RI�鍄x,�2��갾��W��'��-���z7
>��Xqb&ߗ�R ��٣�F�5-�p������AꭖV�]-� G
N(7&Կ�H�|�`�L��q}�ػS�^�����s��6^܏����Ktj�g�ئ]�eF��f�J<��R?v}ߢ|ӟ��M���"��#�N�����+���[����y:�_1y�lÇ�
�vu4Xa�>�|�s�?#���>��&��n�e�F�b3��2�'4�\. �����?X]�mw4��N�'�\$��w��I�_�تZ��aL=���2>��kp���L���,��8r�ݒ�Gz{3Ӷ����(I%�?�E�����!��=uPv�����B�'�Hyyŷ���>W�����y�>N��ۿ\o��#{��]W�c�i��J����?i�ŝ���T���BR'�i��O��}�0��.vʝ`�^��	#޶�d�q-�5�tC����#��*)�{�|Zw����Y�z#@O�qlfz�)�Lk��S�;����lp��Z܎�zzJ��U��Ud��=�M�O:���i�#u,WB��T���d��nf����+���M����#�B1J�aJ��@xO��<���N:�]]��^v���a|ۋA[���̠�T�z��͙d�m�L RcR,,4��f}�vSB�ݽ�Y���t�IQ����z��fF��ґ���i���mi/�p�L©X�JlD�ʤ,�&����ҥ�x�|j��� ��T
>־�@ �8�R#\b�Y�{n����@�����Ec��Pn�Xx%lA&�l�����"���0�/�-��#��|i?۲��#mtغ���#nxM_�m���깮�6��-�a@zH0jcK��#��d���K߽z#�d��������!x"����k�K)�{WI��љ��`��3��k��}z>������=KP��^R�̶Y=ݒ�����#�အ�y�f���|�b�Q"�����c���$Z�|�C��)y�ߌ\�-m�-��'S��4A��R��E L�,pRC�a����b:��m/F���M*������xͽ�78�7f�([)�<Ne .�1_@�B��T`PX�U!+c%��@�	F��quD�`)��Mg��3Ӏ��JϚ5^�뎽�p/�J�Wg8��J��֎#/~�<C�@T�x�e\���A��3w�c�t�;\}���6%�8��ۨw�q󝶸���_�'������,5Z¯xD�q��Hw;Yk��|�vHf�sb��e���rj�����$��|�W4$��W/�(&�?�����>���h��{<w��E7�5vO;y%�/�£���&� W1<���
�R��_}�N��l�@�!d�Ҡ�ꗆE�:-Ur�9c�	Sy�F�٤�&*I·����jIƴ���W4�>��CJ���N�2�T[�˝UYz,`����9cy� @��r��l-��G+����ڪ�s�/�Ő Y �G1,Z9�㣜P��F��p�?�ĸ�mfH�Wj����z��i�5�t�5�)[p���OO���E�D�W��$�x��̢�!T'W{�8��d��aq��oG���U��2��Q�1���9 fy��va�k�����o�� ,YR ;Ǒ�%N�s�Myᒡ�`�-:7��}^��Ш�՘��0��2�!��m�=�7�[`��^<̟j�5�S�N����O����0��|50
L���B�8!����R��}��F��j"��穌�[?t'�Ϫ#���?�Y�q_8TlCם{B͗=��V{y
�7D�������9�r�b��ؔ�M�(ɉ������EVq<��< {�l`��~�m'@�Qp��Z0Ҕ�᪝�:kK�̀�}4J��6��j���@�Ӓ[)؄w��f�E�{��n�� �,E}��Omc(G^E�P�X��A�ݵ�HF��JV"r�e��Y[vS'<�uA3��p#y3�Y�>TN���$�X��n|����>E1p�JWN��?�CG�B���=+^n*0�I[�/)�Y���5��W><sxNI�����~�?�TUE�NyQ*ϰ�̵Fa�\���A���)�C>?wV��YZ����ސ�EX�j��<�RC��Lx��1����zzY�4xz��~�pj^{z2,a�lp��e3A�y�೰g*���BO���4��F��,x�4�91y��^��d=>�5W�XZ'����׭l��g	@Mh���V�:F(�?ј/�O�X�ײ���}ø����ל��8|��:�+ٗJ_��ӻƌ���3yx�	��㸴pɱU�<��������S���o�p"�����{.�+B�/<�m�R��_�'8~k
�U��He-�T(�W2�ɗ��^��(�z�ہ��f�\U4%�jMe������\+��Hx�]=�"�i٫+o��v�Nbq�6Z!��uV)?Y�UΜ�2����!� f"vl ~��TFn��r���V`�W䧏�h1>���4T>�K_����;�2�ddC��lFՆWx�S�f!�f��b{�wW���ko��5�Ad�����W�'>j69 Ku�H:)lIi����G#4A�&��#�3�'�kkX}S�W�"$O�|ni4�NDvD��K���QFPP)�|N/	S�HĒ{�t��A����J䵱�����p^k���ۻi��� ��a�O�_����$m�;���n���:��(mG�6�ܺxԩ�G�;�g-�FƁ����,�m��􏩋�ǈ�0o"�<�Äț��q��p	���8N�B7Ȋ;��*�!-�+�bj��L|3B��؟��ĉQ�B�p�5�*�//�F�J
�Nmow'��9�盝R�?.�(:�&$z;k�����-L�;zA��Q��v��M�b��-y?t���
y�j�}�CWg�Ǆ��?��#�p�K�y�sU�Tr�W�K��	�>H�펝:PkyU��+k�awgf�˖$L@��©t�=���7JŁ��B����l?����B0����@�NN�
��iW�'r%y1ҏt���?hT%�� �7�R�ԑ=��id��-���������'�C��#����y�=|�5ڲ�4�R��!V�bY�es�_�eP5ʑ�22r�P۽�ꉹ8A�x���m�͆%_!5�T0��}�.��un��^��cM≎�#�2/d�Ihր�rf2Ir��B�A���i�}b?�7�;���>���|�<�q��|���PM��87榥�q�mȻܨFTA3�q:����,�A2�����lHS={���p����d�8er�����A�Mv�=K«L��J��h/��I�>n��">��f�T��y8����,�Ĕ@�eJcb ���fti��*iٯ����K�@�3�v!����xy��S�OOO����>%�����IU�ep�'[>X��̱�0�[�iqk��y�� "� �2���I��1��\1���]�Jw�Y�e��M�FM�	xX0�v��@�E�9���<~��%9�L�<%���D~^8~J���a>�����Ԛ�*#c��Q{E���rD�VJW҂_N�"G��TEmgW�E9�)<@@<�F]CC)�M�
9����қ�MI�V�ms5����<lB�Oy�0ab�(�x �{Ϙ�ӧ.)P�fo�W�OP��0��,�����T��+΅�w����4T,�*o6��~�m��,�/��aS��ex>0>W}ܶZ�Ź�f}P��~s�vK�]dY�j�&���hzJ� 8gT�ο�+�m�uP�N`�l��.O�p��4�CT��!d��;6	�:�hZͬ���G��rTar'tC�,��u�T*�j-U���>x�ˠ�
t�K��}�LWQQ�/oW�+�:���OӢQS�^q�B�A��骣J+����GgF� &(]4J��|i��`^�lw�ν��g>�����9��Ҭ��Q����%+A_�*|��4��B�<z�L;���n*~]!ds���ӡ�][��Y�O �*�0\� ��?R|��+(�M����pNҮ'��ۉ���K�!J�5P�e�X���bJkI�p�T5UiB#"P�9��pl}���=+ɘ��;�J��(�ڤ��\!-�kAb'�1̩cH,�,��$����t���@�1�nT��*jו'�_MW�ryTQ�mn�u3=e��.M���k፡��tǽ6�DQ�=��㯝��"V����lx��Rqi��T5���ޤ���h����T,ށl�����JQ��;��;Jf�7�1η��D��z�v��k�?u�.`31�N���?U�q�f�έ<0"�nI���2$�l ��	s[�3SfԫT�{te?���,���$p�6��&sM�����4v���:]P�I(��!��ϓ��N\�|_Ӧ�B�Ӯǅ,�'c�����	Ms� �
�S�(���/#���6�i���J#wb��ŵ�w0�onM�BTv�~u��a;xъS+XFr��J�r�\M-u�&Gȴ�݊��͞�c���~l@p.A�hwb���q�6�u����j�9vEߍ?�i���c��;�V��N����qd�pN��a^����=_! �rE����T�2�oL���d���N;¾'^2�����S��gcb�Y!&a�W��zr�N��+�D�$L��>-�&�=�oq���J�:��������?�!UN���^oI� C���KB�N�ga��ب$Fa�����y$)���9���A�^Zw1���A�
R�UT��r�*p�8A##��VD�b��B�FS�X��)A���P=�dg��!�ʽq���\�)�}ce4v{�Ȩ�:*O��gH8Y�4*)d��d���Ec;_�KGb�Y',YE�67��[l�R�Rk��k��|}_�~���W��suńE��_������W2Mf�'V۶��EO�,b��vС���)59u���d��	Z���>�u{QS�I�5�g�CfF���q����~f� ��f�][����\i��D��9I���g�q-�{0��*t��J
ѯ���?ɦ���>pX<J!�A���z&�Î��$&���G��$Ėa��(B./iP�B��f[���
y��6+C]Ñ|譲��5���g����\�^��G��q���%�����#QF|\d
~�絕ҋ�Ԃ � �"��<�����GX�I{i����@����s�m+���3�*n�B�Fu��H,At�C���H�e���T�,� #(hux��LR�H/�G;|n}�3�֙�}���E�ƍ��(+WB�ہ�!m��<L�Z�.EKKK]0�g�G8e�/~�@��~'��l8&(����%�q7S@bh�zRӎpa�����=��2��
o����*跤	W�*�.^b�h��G�/�!3�g*�8�1Wu|�������S�0��ҍ�+�wJy9A����K�<���rP�2-w��i<	�a��Z�v!jƣ�3�P�}�P��>��W��}?�锚mA��pY�pO��5Z�"�@}4..N��\	�X�y]�ow%�g��.��d��Zג�TP���g6�<n�b��X�C�d��F]ni��Z{�i�K�G#cZ�-����P��\��ϟ�U�\�K���{�롷aU�X/��s�|��T���
Wɗ.��z�@�_3�שF��0��
��b���6r?a�M/8ˈ6��
}x�1 �V����"9�����^Ǉ�ф�$��޴MI���S���W4�dH��dO��{#��ԱG�6��9�N��?.QJ׻X#U����n���ˬ�
bu&���C��4o
Q(�\��h�|���n8�j !�0�f�����c�宕ϋM�4Jo�r�G��j�/�Y��̟i�p;Uɩ�:�d��]ܙU�ǧ��]LBJ5�x�"���_*�u�����f
?67�r����d�!�t)�'�'�-'T<>&q ���
�,�ɕ�/h:���W@��҅0�@�A��k[��˜�lEiP"7��4k�T*���x�3���:Y�Q�!W���c���$����(Fu��eyRtQ�@�ۏ	N���~��|+@��y��g|�� ��E�jg�E��^�xrj�6	F�J.�jA8�-K�Rם ��\���hSմ9T��eK�(bD���V�y��,W�|aMd<�˶s������XP��eT/�Bz�A` `9���Q�p�y�t���ʖ1���pOW�Z�c���k2s�?8m��Cr� l	��ș�`�`Ϟ��.S�����Y#�5�Ţ~��ҽ� P�T򉀗H`?xw�/��arI����?�[�ʡ6���|�h݄�7���)�)��(�F��='��fJ�|��JP�+0�8=�j�������Ƞk�b֌�^D�*�"bw��loΎ"��i�֠`П���q�� �2��g>4"a�È�2䴃�wG5�z�|�����z��N��[>�Ȟ�b�	��*��%􋬉���{��	'�N�U���Fٻ`dْ��)5r�nL�#X��� w f�xS �%��y��6.3�!����<�����h{��\-(��Ϲ|'&.������Y�l�<�Ka�q"����Q;�����t���Y�A��vbW���BxK��~"����!���ɚA��h'��֕}_iV��^�q���l��#@"�R$�q�wZ�pD$����f�8�Tep%`6� ��yA^�"�"v4h��������S^>��h>5���	��J�jS�'���#[6>�0���?�V�~�E�geGd͔hGY�vڦ�deVl��1Zx�vǙ�����z�,�K��$51�Y���v��=�HƵ**�󄫺�|F�:�=_/ή'�@E�*��D���j��vY(�ꚕ���(��Q�,uM*-�Q/=p������zZ�t.�C��|�*�dǾ��*_t�"��֪nAa5�-ŧՅa�筱hd�)�5����ŠP�	�3�M���ew��ˡu��$�Ax��/�?A��~nq�6�و ��0�>U|��#o�왮�y暏���H���V���Y��� �3i���Ж�tY��cG�]F����(��F�X�ߴ��45ZiB��7�&��Ⱦ�Q`5p�S��`%ͥ��ֺ����>K0Pk�{3M�.��(T�71!N��}���\+�5�;��Xc���,�ْw��(�7��k "�p�Ⱥ��{_
�y��� ���7 f`,�m��1��=�}cS���u9�e��A͎J�$8��D�Ư�;����~6�(����
t2@�1=���pb���G����ѱޜR����a��L2�S����h��i%=��y	�nac8�:�`q�Z�B�Yѿ�+9R1	ޢb��|$�)_��痣��Y6o$&�3���J|��L�7�i@2.�v֭���c߁�06&����{�I��O�Q��}�@��Nn`��_�|��h6�*��!2�{`�S1ٗ�@����wd��p4���Wo� J�6�쉌r���\Rr��2���~'yH���B�`ӎP ���%��j{۝1�� 	/!�����(7�%�>�4��~'�ӓ������9��)kU���\g������U���ht��K��h��ޏ���:��qۼ��I,�3����g	;b��FS�A1��kJ�W3�GW���$�9A�1*I�!�TH�-�ђb��a�+#�54�I$���91_N�i�jۈ�U[�Bx%�ֈ׶�������R洕��4G؉�T���t��L�2��SH�* 0M�TW�:^���/�������/���I(F9.�<���"��\|A��<!�"�R?2J�gӫ��'8q��)��I�O�1K�^���R����c�O��c�vd���{e���ih�⾛�?Uқס�p����%�7���*N��,8�z%W��]��m��\-/㲴\V��Y��ˊ_�D�r��赮�%<@��E:�NTt@�&R�5P{L�a�ֵ���ˮ%�veU�&��j {�s����O��v.ƃi�%-Bp��M+�[�R ��ς7Y�J��g���ʃQ6�rX�,]%y\�-�O�i-����7[���=]�Rd(�c�{w���?:�+��g�Z!�rE���G�!�	�hU�$��2�{%=bY��x�~���@�t�ޚ^ij���r�͋�s5��*Dp���[��=�%��b�x	��AS8`^����5��M�1ɟ�U�����:��#��'m�u"ov��RP/o?���GO'9��bl-�� 2p�^��0�W#	}L��8���#jq��^H��Hδ{�a����{e�����P���-$���I�?1o�/�0��֐��j�ކ���������IGgj�Yqƴt�I�F�ޫ)�%�o1��K}���n)��v>�v����;��\|��]�07�|r�D����or���Tv�c
;�a\��mo��.����gn��S֚fd��pc�?4�iú�S�P�Ȓ]�O.��|��Ye�F�o�UM�{
5)���>�E�*r+e#p��?���V� �"`���������>Z�zἫ�b��-Ee)�3��օ� t������X�
�frI�E�5|���-��$Q�����4ljuH�M8"_����t��B�Q�4F�٣"�Q��:�5|Jǜ�{|봌���"c2�{�&���S�F��頴
9�uY�Js��[����>:�Q0/�ZY��;
�N�&�x:yI��ʤ��� V���i[�F�¢D�cm ��F���krFf������q��L_+eW
��E I���igsci�����G�Ά��F)_��?+'��7'��T�Lr���!w�5[
f+[�M�/�A�@;J���6 ���j���+�3Ā��*yj�$�DUeyW z�6���L��	�~��ށ����%
O׷�m �t%X�(�����c�%�~g��r�	q�Fh�/��z��O�t�QR�,��z��j��:�>[]�f�`����!RA�Q��j#eyZuP��t�>-�K�/�+td���-�ͣ�Fe<-�-��A�,rD�FXf��Jܗ�]缛C����������4ܗTF�H� z, �ʀP��ul��TzQ=�����k��B��a�x��J����BZ|���Zz��/3م�9��,]�u�<�3�%���x����˞I��\f�e~B_�.�\��q�2��x�Vm�h���{�o`��&]��O{wd|�k���E榝*��	���:8�mG���%.P�3b��d�E�@YT�	���{*�%���=�7û���z���%��0c���?7.�����Ciu���5�i�N�I���e�d��5<3#zW���ŧ�PDq���I����j�-P�3+�4�����~��9��eֻu�oL�����tt�5��_u
�쟈���)��7�n��u���1���@r\������ŋ]�������|��~��|1ё�h�D�:-Y����E�/���ݶ��t� ��ܘ�z���������G�6�#씍�p�Ѡj�@Y��3����������n������D�ύ(�~'lJd7�nT�w�����}�H9����Jx���H��܊�v�b�MMFM�ߒ��r���-���F��3��^2�
��������!�PT�ʹ}�0�����_(^b�"�$���!��1�{1l�N��L�=nq#I=ʰ�������y�uvꂈƫD�^�u;�F��|=�oG��y�]�6===�@�x�z��G9@��^T�&� &,�7Rmji�x�g����j��������X��Q�zJ7�ȸ3к��/`���좬��ߋq:������nq��z�n[5>d!S�/:��ȱ�� ���n!X�Ť�.�՘T���ϔ�I�Z��#�2�8/ܑ�@��f7�_t�O��YW����ʝ��R���s���5��7����Ȼ#+��?���zMn>�
5���{0S����uj^#��:���#nIy���&���0�����l!i�[89�{q�g��Fߦ����=�N�?M��m�h�G���Ls��6jp�ٔ�|�Y[��%X��6���5'��T�>��"0�G��"|�e���6d�wѿź��/ C��n�?��&t�����@����F͝���A��J� ߯�i7���	:N�/��N蔹��KN�z4Y�!���j(|��<I�"n<c��x(�׵�z��=�q�~�P��G�(5�t���G=�S�,G�u
�m!�3�/�x'ZH3�BQ
�^<?"�0
|w����U�F[�8����Pu�围\~�Ɇ�f�id�j	���i4^�%vϥ.'��3�J�3o�g0b��:V�N��:<���4������/Ψ��C)�39ϋ����p�-���$��)x[��KF��Xw����r~ m7{�`ڽM�G\��p]��)|c����y���*fi�^cӫD�l��Ȏ_�B��J*�K��w�m/P�|+C�\pK:�/��B�l@��t�3��4~�)%!c^]����T��4��&�0�c@g�����GR� ��W�]�b���q��+�H8,)�%���N53��A�8�lU3��F	��=�"� CU�k����BP�`0����;Qv�G��*��a*+��E�F�(��W�s�̠cӏr�3�y�[��/@r�t�;�ۈ�;tn�SR
��eJLN�+)�fM�snãK�՛9�7d�6e&������E!�� �4�Q
q�wN��S�[(Օ���7�DV����O�,*�6A�RX|��J�wr.��0�����f�d6xѨ��*.'玜�a#R�=��M�e�!Ii��ȫJ� �F.5%%����� R�Sk)!,�Z�L�=4�B�Wʩ1���|]SQ!�>==�3uzO\}D�̐>�t��̅p�<�k��ֽ��p#���}SM��o�u_hZ�j=6������G��u�!c�X�x�@l�� 8VV�ݵ��6����1n|v��̇�&��ӯY�qƎcn�&�>7Wy_x^��� ��gd��era8�����2���#\�
R'k��B���"���Q8�V���V A	�H��?K�9��#��8Y��51xI�CM�c�mD謷�����ۿ����v��s]t+�m�g�X��_���?���<��%,y�����!l���&#%%dd��ĺq^:wf�Ə��
��&"e�ۛn�h�얤��*����V.G\e�������E�_��/<a�i��Fmbe̵��ab:��B���8�����b��0�����N����k��.�B4V��F|��؞���(��k��ֱ� �z�z�TF��U�z�V&��=Ø8�� �e;���&.�TZ���_�i���5o�f4�����?`&���j ����Ʋxp\6�L.o�2t�j�����Q��Q�K��66�n#�9C���"�C^ �э�`���|��t����t�˗׷m�;�>�'����7�C��ŏ�F��������/'eK�z�LLL�%AZ::��喔\�0��j�

E�ň4�64&FL^������!((��e��.� 3�\����3�/~N�@��t�>(8ѷ8�� ��9ϢP���:�� ǅtN��/�p2��S70�fl��듥,��A��+��z(AW(_��ڥ����pO��d�Ӹ�w@}=s\�@�RCC�O�y���=�\9r{�xh�Un�å�!W���h����8C$kl���o�d�]nA�[��%�^�]=g�2�bCUFU�)G��+�wG�-���EC#'�L�o�(�X�Q�A��e�?V��S�!Q��%�o+��}4_�ʦ��E��aq��D�/�
�R�Y|�=�{<�\t}zs��P��A|��iu`����ϙ��F�Xh��^]f��6�ݺ�����f!�z!��Z��a0x�W��;�,̸(F�D��M[u�)A�k(CkI	���9͐�f���l%��9
�s�+�ϭ�M�JP&-�I�a���`�J����^
�66�p����.�����n�w�GA8.ʰ���<���d�����  �I������T��HE���>v��=��D)j2�0Ei�8�?�	)$`ے��I����B����ٯͯ��<�25/淺7��`=3UE����4�qR�EOic�Qg~ǡ-@�e��K��x*�.v ���h��r�/��k=���#�Q(�?bK���!E����Ѣ��O������܋���+W�Wv�"��ӹ��/�V�۱_K�n��iT	���f��@�G8rw�c�n����>�b>����{"�ɰΚ�k���-���HH��a-���Gʜ=J5d�a���>�Y��,n��52y�o13|<3;��[βX����A��4%�E&��K���<V(��rScT�#���Z+��=7O!�Ŝ�Z��0�{��&iA�*���M�V�?S�: T{�y�&�/�({>kchM��^RцAH����	Ă�]�BcA(�ŝ㏽�Mм�<r�$��&����w��~�K�ș`�$ڵ�џ/��#��,+ۮ�/�W߬,;'3�ǡ_�8�3W##'�z���p=]6�D�ւ�nj�sI��u\<+�B��� ��7���a�py�9����E�ɻp �����d��}Z����}�muv�/&��S�>�&���nك�iYvq:h���ZuR����H����_��pX:(�^W_{�bweww����s���ɸ�$�`��ܜFX�Q���]Wa�p�
Qsw��^��_L&�Rj���M9yoť�	P-Թ� �>�z�h��
�QQ����T��ٛmA�^�:qO3:q�N��T�m�(�K����H��Ǒ gj������e���4E��-��ǎ�7�s!��䔔��]hdٽ"$��Z|�#����.��`=�{"g0Tu�B[�"Tz�\�R&*x��5��e��W-Ggfjoچ�f��y�@���?8�d�seAi2h�4�{=��k�{���"�p��t0�5��c� s^���u����f�Neҧ��.�_6�"<������5�c��i�7j���2��3> w�?�<ZU]=����g@A����#ӏ޻��f��|iZ�:�[R`Ĕb��J��Ϋ���U#�e�8��,ԕ��zmə�UOO�9cz}Ұ�Q��PR[Rv'����c�C���j�wx�c��ޖA�	��q������&17���+�h&fO�f�Tgk����E��z��c۞c|�M��b`m���K��RK������0�,~p������W!#��+�)�����7G�`"tI�'�agI�
j"]� i:�V��t�6 5v�3�t��ѣ�>O|x���5q�mp>�GO�"�6Ջ�����"�|^
���_޾L��)�+�`��#,?��~�'�PlJ��g�=8�b����/S��a&���)��E��:�����g烌��-��n� ����Mǟz�ERK�^\�4j�=�mO�q"PA	r��>��>��_.U<8�?^��q�����Ç��Tp�@��Ԩyi�?�_�>��K��:X�v�2��Qg�𥞻J| �`���o�z��s܍�w�Z�F��h��L�g�@���lTv9M;�_��F�Y�i`q{�j���;c�ȕ-�y����p�Иa;�̦���p��y=o�{�_�K��/X�V�3�N(�����`�����ah^�dɢέһ�ן�j��3�E8�;t�+1Lf�_|�No��$��y*��E�$�[��fP��o_���}��aza}{:t��p�7wUR���=sv"A	^ɪ'�F+O�JV��Q�%�<��W��h=L�)��i147���2�6�v?0/�@Y	=��_�R�^�ސ��OrH=��Κ�`��md"T��t�W�@G� tbY��l�R|&���5��k��a�:-}�����"�B�v�Ek�n�a�{%�l�X�ݹq�6��FɾAU��HOS�W���i��|�׭I[�� -�U_�(G��2�q��?�;��7�ƍ����������TSK�!�̲A&q�Y�M���C��ZTJM����	]�V�]5��m�ގck치��~��,d��*�H����Ç>a@����T�§��g�3�ȥ��	��'1?Yz+�|����a42��'n��?��VE~�Na�f�+���;{��z|��@-�$NtV����/G��o�ⱞ���o� �Of�د�5J3t���hF;�]�_�<�233o�f��$Q=A͑�~5xhY�N08l�}I*���zsק����c�;��Q�ϳ&�E��H>�!8������.��I�Ux��9�:�h��[2�?�� 06���1� ����0�ɻK�1��-(��<>+E^���P�J��Z}����gZA��}j^�����Df����� ^s�(�C��[���������,��7/bOW�/`�ɕ���Bf�L����,��ێpY���0���>a��)0�_"��u-0���<g'�wW�tY�&�r!�Z���,���h��M=;7��;�@���Q�`�=���o�1�q�4��p���|���KR��5m$봜%x�(bv��+����!q��N�(�f`�J]q��������"5k〙�%*��!��g�Zd�=�]�����;��x�߫��pC��������|��T�����-�T���f7���9����+o�'z�q�i@���M��s���B�+-��:��p����k�`������vta�����;��oK��]~t&{�8�!&�����M� �'/��}�rF�EC~�Znϫ��"?�TH�Q����Xˢ��G�������������9ً�.��6���aeB��C����O ���G�-�W�݌���]�7#�Q��3jai��!����V�Ն.J¶g���G�Q�C����k�]�C;��f���K{�E��x��t,`�8�{��[��������3��E!8�4M���}�ztߠ�x��[̀36� l<�V�3��H�*VB9��շ]��c��yտ�����#@��y*�vY����7�YT<ooe�)Yi��-;���YXО�y���WgIiiO2���
��γ���n���8�ˎG��q� =���#Z2��<xkP\mu��r�+����M�E���!!Ab#�Dq�2JE7�ױ��kR^�#��&7��D7vwΕ`�䫼TcQ�M�Ǡi0�jH�+=4V�G�D(��<��i��@����<�>���2�P��[�lM�_�����E��J	a���1����Wy�t'�Нε�J��4l:~"�h�'޳�(S�CVu}p�"_#I�̾�|l�jt�#�Aa�zz }:Dsp��H�2�)P���Ď�w� x-%Ϭ��i�k"�	��?��
����$�i7�s<ZHX;�s�>�vcsޕ�������)�T"s�",V��~K��*]����Xk��� /�J��.W��,����݅ӫ��~U.|O�:U?]L���98֜�j�X��,����C��;�����o�c��%���2o �U���<��6�V������U�}Ie�,���W+�%43:�	Gɼm�:�` o�M�>��@!^^ �;0ף}-�*9��5*��(H^Q7��S�L�K�ҋ����<�2Ex��п���@�s%��K�_I�c����:ݩ��'�2������[�»�)�9f����&�y�]��g}k�JD#�'B���h�:�`��T^�w4�s
s����ԗ�����.�,<"��.%=��U֠�S�Y�<�(��&ps�=���λ�+�nx�f>�*�8�*�R�Ұ`4�/hߢiQ[n��-56��p���������m����~{��j=�!6�������f�rUZj�6�O�션�{+"�o���@0ˍ�?�P���5�K6w�H�.2�L���I�1s��'2.�H@��Pv�-6���`����ˁɸ3�_��+I�P�u.3!��;^�f����(%�4d:�[:�%1")�6���B��1����{`�{�P��p�Ai�x2m�J�j�"���x���+����AY:�������?̼eP]�-4�����n���]��www�\���\?�������US5]=ӧ�ٺ��szz�F�.<)M��a�K/ ל��rc�?]@SȬ �}���Id0��ʢ�ʂV.�7%�Fw��E~BTn�Ȩe*ur�Z���t=b���5���z!�s���
��9O.yX�_('%�Ml��ʭTt^TgD�k�Hz�Jy����D����f�/�(VC-�X�2�~i�C���%��8����#uw�V,��{޼>`�-�ޥԝ�a*|���ȸbK����#�lB@XYΆ]�y������7w0�c4N�h; ;*	��R��4� &d�#�'Y"�B��.`����R-���3��b��Ä]%3_a���J*_[o4=?�&�(��
��K�������!���F A��A�_W�\��H����<%���z�v�����(#-B#��_��)�ϯ 5v�ΐ���Z(.�'�}=`v�E���� (٥F#���f�Q_[��Sc�ؚ���Q4W�Ȇ�6 �v��:�/(�#�&����j'���B�i��F�*<���"=��>�n�E�dh�ŮdQk.�aN.�KБ��\�����跌��<���K ���"X"â���/�諷��hV�����Zs_,�6}�{�]�-/�!1Xzߕ��p7���2&�LU��)�Iz}Li ��9�4�G��i�2���I�}/���
1p�	�e�5�h�cvL�,�5���C%C^��v��Bf�Ö3OR�e�B�]'x\w���\&��yO����O���hK������zQ$"�n��)�1�3�0\7I}�N����G=�:���T	"m��ϩǾg�֫�W�o���� �(g� �����~��DBb�N��=]�T�3b�����{5{��>T�pЩ:^�E`�T��[%%8@��ޏ����^��F�x�a�ǥ����E�pC9A3r�ea�Lq�O�#E55�`b��U RN_���ū�}�P�c�&^��"�֫���Et:�brig'?s*>&&&�0�P�/���1D
�-�JAp0c%Ko�y��ѯ���L���'n)�v��r�a,b���h�C-@���aH��1��z/�Ŋ�O끁��P۔Җ��ëB]4}Բ'\�KX����Tͧ�ι�i���~�N}V���`lJ��
��ڍ�j쎕sP�#�40���
�a'h������Y�KRNH8��C�v����b[��}"�q�S�%�D}b{��B�U����_��`F"�?=%�zX?��l�U:��I�U'B��ৃE>da!�"�V1�9Å�6m�d�s�a���R"�}A$8��1�u�=M�~��E�	 �~%��R����RE��*�d�Ĳ��Yi(e@�Ӵ�x���t���Uev���jhD�*�<N\��2�z��f�尭̀�ЕwY�j�Q�S�k�,��<)��������!��������c+a��W��0D1�F����M\@�����%�j�&������Q�؜}/�����HD3��F��㬦�J�!���	>�򋧥l�.�i��b[X|�b��e'��E����c,~��ZH����ki�������u]W��N�Rt��!���lm�)��⼥p�/��\	��#���|Y	��ڳ�h������i�ZlRa����c�Rjrs��� &w�kȿS�ςF�~��֏u�t���a�@�C�@�lDM����A��������K�'��?�-��
��{�++A�'��h/$�Yh��a�>4��D�V��������� �*�nc;*eBw-Ri}��d�$�k��G��Ȃe�����X(
LUcg��n�l��>l����w�7�w�<����{<n�<	����}�{#���D�����4���@g��;k�L��t5�p�̟F-ri�xu_��VS�х��k�e2��Kn	4�Ӽ������P-�80d	�A3���i	�������C���(�����%;���'LO���vd68��_loah���Ap�x�t����Op��������Nf�'�n�TS�5�p0��0�hC���`g�̥3�1��s%NN�J�t71		��#�x{�f���9�-�{Z\e�S�L�q�)��3��-R��
��K����:-cn��������RM=�m�*�թ�șl����s�@�b9p�ŗ���:8a��'xb�g���h�H��&�����j�����������-om�ن�IB��W¦�>$����F	^�Q���MC2�!�Ũ���N� �ћk�$k5��1��F�7�=�.�Z�K~p`���F�Gj����9�6u84t?���Ox\�`��M9��H���Yg��}j\c�'Rk�6�������!��W>䕿/��5eF���pTS�94i����:%�P�/�\��}?H;@qi�3�Y*�~�B� �\���yW�g��G[����*w���b�.ŗ�;�؟��o��ˮ����\o��<���Nw����v���Д���k�m����ھ|�� ���9�������,@h�#l�~\�j��G���Eڲ\?,E�	g�z���j�,CU��c��v__�wi��*���_ؕ�����M��B�;�0wV��#����)a�i��}P�q�^�;�*09��|����Q5;�9���y�K��B�zW�E/�>��K���e�Y��Nʥ�hggGMO�����k�=��k2-�{_NT���vMy�����kZ.�ҩ`q4k�8c����)�ZB��S��w���8Xb���[:����u �L�Tuz��ɸ�SK�*V7nhte�BS�%%M-�^3�V���5ۨ$A�X��&O7G}g33��E�}��222?���P.0U����Y�T�K�� >3�u��c$��-��T+j����\�1��La�-͜���������%S��s���LE�;}���:�t6�&�`�4�{�$�s'���s0G)t���Ů�%>������v7��;�	�+nzv�J���m��-=��()99Lp�� �,��(e��P�!����,��A'�0U��k�k�nK�B�d��{K��D\����C�����3YY�@(45���vg�!dl�,K����`:4;�ڵU#vq�d�/�� 팱�ፅG�#b�h�I\���N.S��B�^�#��ls��i+��a����wr�T
ף��us!�j�����P������<l㋍M%�����7��[iؙl=M�-��� r����|��v����H�?�~ZML�&tZ;�[ά/QL1`�.�>�V�ٹ�jui��۱��5���^�Ze����S�l��#z���𘹑�:c��)���29�?�Ά+^��X���"�2Y�)x"��޺���������{b�����f��)�@P>���9�A��7s(���Q��[X�o�s{s�"�Vn�:MI�W�m`i?�!yq�x5�צ6�茥�_lS"B�sr��+"0�4�Z��}ó�'y�1v��k������o�p�\��rI�H�z�etY�ۻC�U�7�䓍�SP���V#%��zT�4�M@�8_q6�+��j�Ǜ}:D/|�K���l+�"�!)%���ibb�^xz�5����'7X���'��6�E�_���9��u�Z���5����wD�,\�BK��z�+���;bv{��@��	�e�Xe��'�ѡ�ŝdR�}@�ߌ�k�Ғ�m�6"]�5�p{�hm\eaf���W<kyr����dG�����yL�=�j�`�����V�`tO��={C��f2�(��a,�b~0��;��w	u�wk�ԍ$i$��$eL2�2�}]h����i���G{7��x��c-�yFi���aRE+�$=��W���+��-K�t:b_L��ʁ))��p�h�b�8͎���dՋ�b~y���&	������-�{��4��Ѧ����ͽkTw�p�,6�+���aB��fλ��-�:�8�i�+:�7(�%2���L���:�����sq�M6� 	�-��K/����w����ְ<�{5Za]�L��Ĩ4��ˊ7HM�8L��0h����-�y�}�l�hD.Սb*`@R�B�]�.���j�yu"Q�X��RX���f��A�ʹ����.ռ1����:3��a��:V��trq�I"؇��o`;�%�ٴN"w�� V'���[�R�f���kH��sï�FH%6��9�"�L�Ͷ���$^���{�� �A8P�AS�f����v���czv�d.�H��|�c��r�]݈�j3���9�1z}q�)�Ml��=�����kA[���f��F(���������+ZN������4D׸��e|0�]02,v��f���*��v�~��|�,�WrAA�o�%*��wR�+�e��k*���s�F2W��db�Na����"bSJ����n��Ϛ$���~a�X���{]l�'�;��#�2����T`��mi���<~����F�)��X[��Y�:d�Ȱ'��A��^�Q�Z�i�101�A7A���D�X��
��v���,=�7gQ��4k����<��Mz�I��Q��(��j;���WĐ�T������V���w,̕�tΑ�T��x�&��/�>%G���YE�g�n�_�N ��u�)ǝ��-�J�!7WDP�H:�!m��C/�Aۨ����mN��qBp0�\���a��C��H�2��c��������X8!JÊJ�P���W��֤��J�hS�]9�12 ����PŨc��S�O�)� I}Y�T;4Rk��'4^ʶ�a�vǧe,n�ժL�L���θ��:���mEi�G�3��_2F b�7��C���E�����6#l�\e�TSΰ�d`������) Cp�Գ���=.Fp���zI�.�]��<Κ�@J9i8/~��������5�풲ʒ\MWf^�X��c~ױ����� ����+���`ӵ#�C� ��L ���Gh��X�pz膤�"3�������*�)���Țg�/�&�R��&-��0��$�;(AT�����!��x�%e,|�C ϶qn���.�:�!=�oz{{;�ɜ����7��I37{�j8,=t����,t�
��	<��n=�:�4D��j�H�k?�G�&�<���-aqB��g��\w��&
�֮F��N�D��h	�/e1�����Ke���؊�{<���eH�T1Ě�ZK"�i���W
jЯz��eP��/����-����o��{�&e��Az�X���N�~����Q�o\�2w%�P���È��,��*�b_Lx&	�a�9T�v8ߓ]e#c0�P��0�Ӷ��s ���޴ST�y�f��xD~F/��Bbjj�N��}�U����E8ѭ��7Gs�u?����8v��XxX�l,�z��D��}�vF6Ч���9����G#a�_�/���_] [��Wd�c}x�8=�V,ϳ�x��TmaZ���ʵTȄi���(�X�8y����a��^g3+ �BEo4f�Jp�H���Wb$��I([����Ԓ�ꡏ��߰�Ο�t����g� � c6r�/�=Ruba��!G_����rb���$��q�I���F�����7�Ks�𒓓��PlͬhN#h�&�X �t��/ߘ
J�3�����χ*�IŪ��QI� �����Ju��90(�͝��*@f��1�+�Xp��L����� �#n�eDUX�f���qu���|M��c��b�:��U���]���+��*W��@�EM7�3n���4����7_����3d��b$��!���Ґo���{��A���I�9s��Z&C���Jq�����+Ӟ��%!J��վ�!�jܮ����莾��4��:#�"������V\tGc�|�9��w������v�J�Sa��$����9�Q��3(��蘓d�7��k���+�>҅'���O|!R��E�(�Lf�O
v��}D�xz�x<4p}*�g� ����}5�r��
Y�g;�)�*�=��`������kﻘ�N�;?�S��X���J|
����/����x2�,V�@DP�W�q���mg�����1S�`��3�:��cpt~��:���4W�R���<�;��W��'�n����?�RQI�a(��$�S�@���@@��w׼ꈽ�T"�E�j�xk$��Ţ?q�q�C����Z~����a�AZ�y�����@����5�ޜD�T�^/����%=���F��(g��Q�mKE~U^i�=j���p��k��y*E.r1r�Um��� ��U�8�=V�$��#������U��4 {��2��jGS�A�#���p�H漣�����q7ʨ%�.>��/���7��eSQV��E޺&^i�D�˸��t [�#"}��ދ�GR�'�1@@/�*�0�8�� �^Y���y�d���Jc"��ί�n����ۊL8�S�i���t)�?8�L`3c���h�����"��hu�$`�zgfF���a�H��c���J�Z��1YG���	�x�=z��˒c���Y�`2�T�ӒW��A;;)�e�OGLD�,=������O�R�no��$�������)�-�jd6,�7���������{4��d>��䐊1/!۞�4���}ϻ/���X�2&���|ǃԍ�������W���}���?Ƽ�h�����TSc(5~T�	J�#u��Ȏ�D�ImJ�)���V�@�Vc�p��@�UD�r���վ+�RR�Iל��{�������0#��[�nX]	��/�|v�h6��ҶK�F������vH��s�|����_�2J�Gqzz:,�8./���"B}��^��7��I�̛���"�pKNO�����7Bǰ?yo���7+���Q�A��m?�o��Y
�+�|W�xB(*�©�ՒJgGTb��0p�]tc����Q��̂V�L�R��^�w[��a �R�@y�2���8��D�ܤ��$�Y�2��UԼ��	.^�BAS��o����`=������J��r���������0�:��~�B"�l��ͧŖ��H&�92� ~���#��m���#���m�<#^�u�L�r���5�FH�'����*�?�	t���j�ށn-A��֔�7�I�]�(&K����O�jT�XTjo�������y��$$�Y|�k�z�멜�� ��J�KB�Q: 3��J.g�b�qX$O1��Wg�vV�`�)i���ҏ����3%9���C��-��0q���vF���1\�^�p���_���m�^/���i��y��0�ԛ�mmZ����LǷ����}��z?XޘV�wdMmT�Uh�t+W�V~a:a�j
19;;B|LxXT��eYA�R:����Tt�By��Z�*�Q{�rT;�Ƽ>��\����� �D�>7w?��
U�M������^ތ(�쾔�ؗ1e&XZgs���3�Z��jun��
|�B�xy4F���@�%շV%X����bhy ���=_ӫ=[B�^<à��5:)��	�~� �/�z>�hcg��WXX(
�����9�]��@r����y�a�T�AJ�}�9����6�� �tܾO�)Q,�6�(h�ufQ�bHS�"4���aY�`�{R����ښ(�����i��-ˇH676}k�+�>�_q����]�8m�*>]sI{dY]�IC���u���� �gb�@zn[�9"rr�0�h�ۻ\�����.i�8����d:��EL2��֐H7\?�)���ӫx�\�5�U�,�����\�PCII�;��S,ӡy��(��JG�F�����v��Ugu=H9��j&����U}��gF�;	3�B�vj�0?��iww7���oG��j����xg(�9 ,&�H�(�D��ħm�:�R��~����&�����N"��#�F�2�`��Fv��b-��3�oNu�i�}cC��B��aTl�&��%���8t��Н�I�DQy���GTħb�&�^]̲Ա���333}ώ�g-&d"��O�d����a�h�7��3S�*�����+q�.D`��O��.0�>�+����3G�L�1��օ��/�N��6�l��ŷ'��a�
�,�����0+.��D-��[�����j <BリS۾��472I)K|�>7!��4&s�	�/���t���.���!p��c�B���z�7]�JMO���l z*�Kn�l��$�I�����G��ő܉��s�d� 1�6F�t�V,�]�ь	 I�'4fp��՞9c�Kz�t�i�����"�e��unw]Tw��q���`'^�O�)�[�=����:Ȝe\S<0�stG�8�VQ���J>�G�h�ׇK�x�8a�^a!302�H�'i#�>��ྮ�\F<XeOC/X\؜����o�NԂV����R����~�q���ŕ���л�i��-!�(�r�c�a_ey������W@յ������+��Pϐ�Ɵz�3[�|��Yps޾��ʗw�x���Mľj���~�Z���&�t��"�T.X(�ȍ�>M""P�5��I�S����x�%	��ib�:	��Aw�q���h���F���:��ೌ��b>kl�j��tm1�v*��C�U���^���G�'I4��1���t�d�հ�=��[q�j���ʜ�z��+���؉���Yb�P'��[(���h����%��O>�,'C虥��0<��sǈI�Dx( ��E���� =	7���R 1��(:��f���,o�F�_�O<D�P������݋��]�� ��ը���_�̇��b\ŝ�0љ�u���EL�e1�9�4��~�1�I�ݩ��%�cNO�%����
��9t�s�$5�!!%?�bF��,�B�`+��b�H*q-�7[K,������QX�w��86k
����]Ƥ���fie��	8& sP�����3��-��I[���+^���SC"�օVRO5ǽ���8��w�� ��$Cǜ�Ѽ�����9A���bc�@HhOVn��4�о��0����]�V��gR�<��0��2�'?j*M��p�T�ʏ�'��YG-sNb���|�.R�����Z�(��.�e�,q���$;����ds]��]򲾐2����:��!.e�1
om)־{A�0a�`�k� ���ފM����<1�#{9�ˬ�X��Zm�`�������q�`i�g�M���-��q�%����C��&��t��&�n�AF�hT֙���|����d,��	���4r��, }I�Fj��;vB�
>[ô���s�fY�#���E��f��3�����`�q��O��:�Ȅ:��[��݅��i�ǣLts��C���?����:������)"}�:y����j��X�r�����O8�EEQ͸������7�2�)䔡��|v�4��!�]n�F�z�*,��a��n�X3z��-������ch�Wq�沄����<o�,�q�ߙ/���;���>�5�������qC��O���b�!y��K��45a��~���"��Ǐ�gWy���b��1 �_�&�t�2?F��i�����v���a(��گ*UN�pG�����C��>�,�_C���U�_]�H�b�1�߉�v������X������A��	��+
�k}ݲ։�U����{��l#�!��d��3����1d�'��҅p��7��/��!�S�G1�(�V������bɠ�H�8��*���x����	gx�+�%����0AD�+�'�[]�Rm�JE���t���4���=%�X�8@m���VN��Yu��C�m7|R������Y�O=]5X�*��� _Ո�	u�-^ǋ�N��J�$�J��� q��(>�k; ��(vO=��sz������^�d� ��T��LƟ.���o�L�k������B�j�C���Օ�ʔ��`�HX��K6簏�l�³��/�����P$ �Q��gXs�mWy�p���an��{6�	$���J'��P�t�D�	f�pk�d
���!yZ�ǀ�+�ޮ�J��Vǡ/��/�G�.I2��Ƈ�nJ��N��jWgA
|ƵM�Ex�d`T�#fM��t���{r�<��$)��"�Mia>���Ƒ�,���$�}m _E�yn�o -I�Ut��va��Hx$��)���JH2�m���:�4�Y���(�L_?�`3іL,@�:y`�g�ͷ�Gi��3���z�џ>�[��-�/�^A7����������"���-b�d�m�����w�>�Ҫ�w\g��ܶ^������HR��{�r�Ff��Z:�#�^�N�
w�jb�\�dBm����9E��o����L��
S���2 �$�VC�n��<����%TȊ�~v���@���Cű�
���?M9���$���`l�`\i��Pv\���� +�Wj;3��y�<��<U����aC��C�z��P"��R�
����/��c(V� ��(��7�Ǐ�K�NkU�ަ��P_���3��o1m��}�jxf+��M��s<�i�tt?#,�s._6�)'M��I��L\�:�őC����4v�4F��	�Q�sZ��Y��ۅ�_�=�9�9(�	��E5J�(DtS0\2P�P'�Md�/���\�OP6mj��ʄ:�`<�X�z�'R��э35�)�U�⩹�jNv)`��/�y�\�{���6mM5/�b�@��^�.�	lܾ�9�l���\\� �Ux�,dם+oa���H&�1��WꭴA�%�Ř���b�S�oǺ&���J"�;b��h��+1/ 0�J��GqfB����RM���!�˘��m��x���J��$��ZΥ㢶>�@�1�	R	y�&BGĞY����m��8� �D?,R?L7�����"�,:�(�F��9ܸ-���7�|����Y�p�ߞКe�:,��_�!Q�H�~����Afb�%D5��_H��,�ϖK��WkQ���fG%a�,�ef�Q�����d5A�^<���Q����ԥȊ�	C��X.���I�Q�
\ΤH�L���Ф�2�ʸǩ��e�_3��To�&�[9��jة��xH���h��P{4��~glv��r�ƛ�ܞ,٫�%k<���0Jvf��>�[��o,�"Q��ڶ�����*�H�	�kP��0 ���2�K����BRŞŝ*����$��J���������9� �ە��Q��\"c���"����>��'����+��xe���ŵ�҇��QM�p�6��!Ǵ@*W/⠧]"���'֔�h(���ֿ@�f��`���`j�%g��/8�:�^m�嗟��B&��[q6����5q��z��!��*��<�z=߿{=).s����P�S��<ʗ�O�<7(��/�)x ��m���\ ��k���4hݯi_7�yW#�j���6��R��C%��M��xO�$Ә��q[�������V��v�
����N�l!��Ls���RZˮ����W\���Ze��[%�3%']u���Ԧ�xz}�g�¨�=���`���}x%��p|J�(��.n-���{���^~W1��+��iQ;K0>���s��ye#]1�����)����4��90d�\����pNr4�yw��Ѿ�]o�k�d�
���m��_�?`:_.,��h��	���u;I	*��k>��΢*��B�F��S�7�q6 T�>c7�R���K|�/��sU�����$i[������o������jϝ���Y]��Sg�³�_������C�W�	�㌏r<؆��UF�<� ��v�r�e�����W�>�:_�yꮎ}��l"���Q��aD�BԞĦ��y��N�=���7��+��:�|/���8� ��{���LJ���g�9�:�g��b��RbNڛ�O��TK��F�F�+5��׳Y����qT�Ԥ	)Za�OkW+�=��	T�|�\�(��m=����hM��Bz�yb���"�w��2rc4�|��sﴙ��V`Dz/�.�qA�/�Q���+�̼�P��=*�(0+�-O�+�%����n����b������ԁe�E�e_U�Qp���јZ��rL��/���8����`�]a����P�H��ɳ���"ȗ���+SWs�}�i���sǥmٖ���=���:���+�!���nv���*�f����ԟ޼{�6�>{D�imR�1~n[=nG�̥W�/�/֣)��<3T�G���$�0I#� �'��pE��ki��r\(��.��{�<K!UD[?S:A���{V/q_ӑ����gI�~Ji%�WMJ������:��	�1|�А�Z��l���P�ǵ��Qᵦ<S\ퟓsq�>��K����X+�m�Τ=��.A������)?������L��.Ы�`h���q�)-vHf�lg�Z���1"+N��������ف��Iͧp����L���E"��6F�ҰoZv��oJ��QL��J�n�v��{o���bkݚ����� �>����G�ҝRW��a(T(����405�V��qXZ�)�S�2ͥ,B�L��Ha|����Z�gٸr�H�/���8�Vӎ/���lacs�L����s�{�ړ[����ࠫ�[������:ź��I�-ʽOߍ��%�s��@�SW΁�`oG�n�钨(��k�#�G���U��`8�`�jx��r<Ý���&�`)۴ <t���,ŉO��E�=�jd}b}��|�d	˥����G_�9O$��nE��dH;�<�_s���X��	������)�����)l���ja���QP�HT�Ą���K|4�y_'���e3�����B^48P"x�b�twmYu��W�{n:��z��3«/q�W��W���^u��y��devg��-��+2A��nw'�l�i��A��@�J�/�Y��s�AIյA�(��r�7R�9�_�#u�E|�vZ=�S��ݘ��!Y����z�S�=�kL�Xy�Lawq��a�>���;���I@���o��R�?�7�,8�,m��1�x���<�A@��_vLk'!��ԈcPMf�CB�u�S����@ۜwW�};`qFz^U�.8���7�����&I<��ٰ�Kx�����?�,~5X�w��q���b�z�W��z%mЮ�>Ȋ"-§0ߋ,U�L%��>l�nӲj˙���Uze=�d-Y&�όQ�h,������ 
mgQ�S>ە��voӯW�jsu)��`C366�K�F�i��:��х:��ک�Pvn�Mͅ��roP��$ ˀ���!�3�1D�p�߯W%�,���T���;$��7�=�UL�HU�æO�G��i�4lZ��:��Mk��EI��Wsx[�S�F����+ʿ��
^[6|�N�4ʥ���1�͊Lj�'Q��d �~-�!*�-XA�E�N�`	$�_\Q�:�z���Jx�u�*��'n��7HaJ}��D���Katq!xe�5��!:wgi���kߦ$�=/)*�,'|]&�;�%}�I4o�t������*�.rv�$�PcK(� e�i~&�V���\(~�f�ZP���|���Æ�S��}}U�JZ����#OG���Β���DA�k�Vj\��5\�h0(aSҪ
4�����@!w��~�;A��MOZ3�M�&5`O!�������Dά����1m����d-KEy@�_0܊,v1lG�J�`�T����?�G�������/mHM[5 9:[�%9&��?u᧚�	=��w2�@�t�aʰy;ɖ*��"��l�u��עs.-���ߓ���Ҡ�]	L�M�S̐1�Z`zc�<R�|���Nz�/�J�2[���)@t���<(h���|�RC#Q�Q�=I��� x������О�
�{��!z��.��[�������z,�é�}��YT:C6u �p )�ϓ�y	`%?��T��\�Py�3�b��m`5:����@W�����O��nH=�v)���N�Ɨ�\;��6�p&�8{�u��Β����+�i�E��g;%.�r��;XC�}{�� �ɞB#l����� S&)咂�����j�mH]�~������e��'��|�6WK*V��٦�3����j�pR��%c�R3��c��������ƯD��b�	Q�h]BԸTi�Q���K!���r�;{K͖������dlCbt�w�wu���dxB�ZU�C�0u�`�NLX�q�3KU�JJ�@"�/E�胃��ꉣ݈g��s̙v�&�:��94��r�>'2�W�_PM8#jh�z���_\vv�>�����I�@U"�>Bx�L��Y�F#��4`2E�OpS2�\����j8��d%�:z�3�QC���0D�p�bWBƖ�A��ՙy+q�����5M��H�.���^]�r4����q��ӉF]էit�b��V3e�p��R�tE���,&��
�܈�Eǭ��Z�yC��}t~	���\�R�� ���
/����hq35�a�?��q2m��}Z��ܨ67�4�D�[�1HѰ75�j��+l�ڪ'�@��t�+����-��},w��ܘ��%�#@9�fxkb����ih���,�4$��#S���������Ueճf�*/�u ���]�=��1'��<w�C�{v$@
���rY�� @ �TZ_�ѝl,��xG�e�%���{���!C�lך=�&�7s��㓁�}ס����.�>�6�8��ƃ��6�����@��4Ҩ����B�>�T�g�w\�@\�F�yL߇�U~�M`g���ڬ��ݧ��!n�Cq�_ɝ�����QXq\ 'Q�YFJQB�U#�u$n���1��a6��5�gB<tvT�f����FX�E�4��>޳1^�U�߸�J�q�&�U_�����'�,x�g��yHw��X|���͋��iҥb�.�"Gz6�	S�4z��M���������^p�g����Q��	�6�{[�r�t �m@�釭�G9S���;D�r�	�M�uC�'S	�FB`��v7�����i}y��܏��c��{�>�����v��}��׆ݜ�Դ,��?f� _�ˇ�e�0�ȃ	;�}�/f�����?��4G~�������#1@��;�~K�W�����B��A�v��苮n̏�]�e�$������[xt����h�%'@>mʽ�y.5�H�a5���7���O�CӶ�%�5wj2`'U�N�H�	�P�(����7����	���OVN4�w�ɂ8m#���L0�J�����ͽţ7	D���75dW��E���ߝ@���m��όuH������"	I�l w7-ll�á�Yeo�$h��S>��6?N��0�xԩs&8��o�Uq3�:���1���� ��2TXS����sj�~axR� q���[�����P5ŷ����=�RAj���u��~�l+�P�9xVU�,�Y�i�h*f��l���އA��-�&�#�k~Mx�A�E��ؕ�I��RW�϶��s_P�w\_+���U��𤣓��+%z�	�9�~�b�����]�<�Y����R�<Hy�s4@0g_�i�t�(���XY�zC.}�r�B����}����/��ő)AR���[U�H�j���Jhh�R�U����5����ݕ�%��Nn�xD�6��[���i�K����Ga�Q���=��~Woy�l{ٱD��[�/:��ήE�J�nܜ���g���{��b��Ef�f![ $̂j�of2�o|�Mmh�V��d49�i�$��q�����9�Y-6��咒EWy+/�>"*�r7��R������(<�m�є<еM����D��T�Bu=^g��>�W�ݒ���$���8/	��a�5��;��(�~�Q��8��.���P��9`��J�����EK��0e�Wffv�,�R~��JLT!�%4�7�̌ɿy����6R��c��S,g	���d�����W隺o5V:b�}3���6rmkhK���/H%�T�qe�1g�=�9�Ő��)��k�V��Z\�WO�JmW2l��O�4�)/�ݼ�)�$ѐgHE����1�kO���W�抿9-,e)�d�������.�Zq�te�J��m>whՈF� �E��h43VC9ǜ�3͔\�b;�7�9�NG�t�bhmnZa�Jy��Z䵵5Tt��
&��*U��T1��J��U�cQ�G6�3e*vt3�DŤ}�����i($���K�G�#\ӄ���c�r�\Hɓs����
;!����������	��w��.���E�1Ŀĵ�=�:Q[n�|P�ҝ{��?&|�+�?ư�	���SH9Iu�A�nn���|���T�Rb�O
:֢3"��D�� f ���Z�,B}�]UHga�j������0R(��Ae��p��ϩ�W��=C�9��a�83ĵ+]>�X�LD��a�9��i�/�7�=\7��IٸH���=�%"uBӘ��~��	 P0n��3_�7�}�Bqiqw���Zܽ�����Cqw��@qgp-�n�=����O^�JΕ����k��dFp�XfddD��]M���t�7]h��Ҍ������B�x"	��Cq)�D$e�@}
�gA�Pe��_i��t���*)#�2q�݅�^��.{=_���O�Ff��������ϫ�a���p%wʇ�\�	-�$FW�H�H:T��m;�D��H6Y'�~�s�l���>xݲ���H?��	,�pmxܤ�ש���Ef�����u��+-�<�"�o>�}�[M�"��o��J��0{�<|��R;1�hz�% q;��2BS�,��]�j�#L�8�r<XpӋ_�=e�s���ޔ��{)��ڊΫ���SuJ���#B�<)������@z�Q�I4i1��c������<��Zq���6�Z���޻������}Y�Z�!��+��WkT�à:�����(�И�����Yh����9X��)�{q����G�7��xæp���a7׳�:�����&�3&����S�m��|��
�Qr���ت��Д��	�}�ӧ���D��r���ܖ�-�ڈ�*0�ܭ�ƨ�p@9�rw��pD�����9*��^�[��O����X~F
97b��<��2<ײpss���_�kf'TS��H�e��G�x���}�{�x�Z��{�0ϻ� ��HW�/�	jX}a�ٻuk��$�/�W�i=�9�+f���"��ҵ�AT���.�VV��hoO���}
���T��1kY�^�w����|�8o�0"rRRRr���vW}$���iM�%б�g�_�����j�ƹ��e��z�;M���/ٲ���t9q���2��Dk�ޛ�Z�2������X�3��jS�zU�NY�ˁm,�����L�Yl�����"m.[�tDd�JS�4��uK<�hɺZOrb�Ϸ�1R�Rc,���̊���Ԭ}|R�3<#������g�ȝ����q�x�).��([����",����ٶ��Z<�Z.ؤ��삒qm���v.F�E�]���rj~)�k��O�F�χ�V]��q�����?ֲi�zρs��0��vj�W�SP[��ۚ1�{��%F��au��&!��9O��j���JV5t�(�
�mi�]v;�K�l�je����ZK���.�VWNS�s��Y�S��+�_��;��.��gq��\v�z�~�o��%!��g=ߔxY��2m�&�R\|e��7�f��3X>�
N>��uQJ�ð����C��U%V�^��׫����R(q;zLqI��)P�p���>3r�J�	�id��r/rϳ�\J(��A�1�v{.���	�%�/g=�b�o%�veHG"b�/;D��5&wg����q3b�)�v
�G���t%��gzy���Sh����<�I{'c���a%����x����f5��I*)��U�T�{���B�F򙗖��c��2$�6p�6A��o4�ʯ���@k	�<\1�&L�F��7��֨��X���٦�,7"�n��kmB�Q8{�ҝu?S����LkCV$�78�O'ԙ*2u�p���I�Uй�7�d�͹v�포R�����X�o��˧"N_�=�2=��֪_X6dD��n�'2ܡl�QnF��!+�@J���g�Rqw]ܽ�Xry|AUv{�8r�yYiOm����W��x���~�/ګ�}�,�Nt��5�@�_Ț��/m�y�o�2�3]��WV����w�[�ꂀn��p��"{I�|N���%�$�d��}� �$������yIΊԺ;������q�{��<g�Y��߈O<��n勭hZ"�j�Y�K�UZ�)�(�"�\=�+�e�"��GD0�_�E�ߣ ��^�Ɠk1�Y���ɗ�興j4�7(�%�{ZWӝM�s��ױZ+��� ��\®�Y5��[�����m�z��b����L�Y�׈>˵J�qv���j�rWM��W��xf�[�O��H�b2�v(1���e)��._N����Y�C��s*��m�R�%Z����5!_�|6UCPT�qX�HH4aރ�|��JW���#ܹ��^��3P��n���K����kB���}.��f�΂,���������H��Ŷ�@�A�S���X��t|�ER/V<�s[x�4�:nu#|���85cv`Ԩ,�<s҄l0T�����.�S7�ч�@I��S��2�żs(g��b��4 �lH?#+��@|W)X��4z��W�;*�oC �Pv��ߜ��o��y���5Ͼ�/�h��רI�04q��,���G_���n
p���9/K�66�\q���yA�&̖��Z��<��[h�<�/B��._��<k[��w5&���J='��ۨ+NvҔ}*��mJ�D����A�E�j(�P$$�3��݋�����?�cs���L��"+��^�[-���kM=&���?ɹ�H�-{�[�����׏L~MJ\�@]S��X��T��\�a���&���j+x+Cɲ����Zޖ��5ed^�l�>�pDrJ�h��������IԂ:�(��Oe��~�+�F����F�����E[[��?��+O�C�2:,{w�2��d -��z��ǳ��.��X�����n��x%ˊ�� ^� ��GI���1]y���3��+OoǿW/\�.d7�e�~�c�k��c4���Y�:�q���|����WJ�\�Ȉ��[����X��OW-�)�ax�S/7�ĕ��wS} U'�,G���}��P�8a�r�ǥ5Wi@�yj�/^�͕���!������p�/r�VO4����>������
I���0����ěN=N�n�}�(��ў��,��L��7��<�������@:�ɠ�ne����T�.@�����h�ͽ��BL����t�o�1[o�4Q	�٨P�P	K�Y�E�OA=�s"t��j�<�a�jbbf�]�+��Yt����;��ӧw?ST�0j��a2�+Ύ�l;�e�L�sU�:.�|����Kt&����vTx��U�y�����8N��i�_��3�sS���ք��H�x�,�c��0�tWc|f��ǃ�z���;��U�[��28����c��<F�4��.����}�Xi:�E!�G�9m[��g�����i����T�+�67����u��?��·�P��q�X�s�\�!gƎ������������h�����B"?�C5����șR<��� ��@Ўvص��ڱURђ�]�%E؆F���Ɵ�\����-v�z���/�i�v�����M}v����e��khҝ��� r�ۯ���D�"jᓒ�ͽ�!��/ǩ$�������<uu����æ|�g3å�d�>��w'�6c��.(]<}��ut��-/RR]�oU3�Z�F3y�9i�/����.eP;,ꤾ;f�"�0c
y����,5=J{�Ģ�н��ֻ�^�����3h@���k�_�9����ȋ沈�
v|}���5=+�dup�s/	�䄶'�;Cq�<�"�w�g@��A~ϳgL˳YOYKr�Z�������i�k�����)~Y3��ǻ��"@�p�)�*X򒲦ݵ����`��Uё~�4�͊Oϑ�#��H�'�������\���oЕ�םg���=��;;r%��=9|;��p����6k�2^ږ8��
�125�ȫC�Ӥ�A��~s�̾?�9�\���9yo��"iI�"$�F�J�[A��M)tk��7�s�
����@��/��Ƶ���A ��������n��^����lQs��:q�)f~�W�����p�[��Ew�c\�j���u!TM�1;����{!3^���{�R�]��2��E �p�r�+��Să~G_��I��ug�Ob��}2>PG��rڛ��6�?>Q�k�9�.� O�/�ɳ��c�@C�K����3�:�.�ܓ�@�u����/ĸ�Ʀ�ً�d[s�c���ԍO���Ρ�U|M�q�U��bYd�4}������|{0���Oo�n/�4~8��z��H�3)�{i�6�I0a���V�x�6�����[NuI�	��F�U���+�	�q��Ԕ?'$j�r��n_�&16M��
AY�,̕*�a��
�N=B�[��x�F^���	z�/�OL"\�2�A����S�J��>Mݿ3��j>Ɋ�lM�S�����vS��:��,��$��H�LH���_��u�X��N��s~rSv#�?�Y��mCHP_������ΐB�b�Ό��矬�ZU&��h8��'��5��\�+=G:�yl�Y����+>��}@�����4[�V�$�/h���!D���#�
��e|����d <�$$���% M���7��pa���Y���T�JTRҨ�/����g�7�%滏� � g���]��ߵM��o4��щ����I��F�!C""b���o��~)�^�[}	Ҁ<�^G�=3�f ���	r�,{���i�S���(ю�T�@j�OMkՌ����5y%����?/Ǩ&-4]}�,]�(o�þ`�hk������̺=�;�`�9G��:����y��UPk��)�s���>&Mr�ٷ��s��0�L�(�����A5R��B&W��^,ӳ�����sh48W�U=�&.U����7�/���%~?�Č#T�w�SƧ�Wu�x/���um���}^r�����j*��©�aux�P���dҀ��nʹ��PF.�Z1�� -�߉��&?��9�i�(H�������j�O��ѩ�UT��j�{ڠ��	F�z8�lo]��6�Y0MѨw�qL��030��	��Ĥ�T��0%�t�7���:��BJ*C
��ߥ�)���:�7$0����	�s�.�FPA���:�eǉ�&@��r�7���A��K����>���X�FZG��?���%0)�O��2�IA���j12�~+7��*'�u��j�Q\��ed۱�_��ZЈ��=��zqm*�5����sJx}X7�!��w@&��Y{�����쯦I��B4����y��Q��0�_���[�|��I#I�������k=[�s����������=���:n4�C�UIԨ��v�����{k���.|lu19��S���^8��;O�N�4梱q<�t� �a��#qc��{��}�gc!�w0�v���\8�d�Q ���D���4�yF�����V.u�׵T�}�0C��G,&����O�A���:]���{������� qB���<U�f4)�ڔ��?�%����<2��8e�"jȣ嬄�8���AF�g�e�|�~�z����!��s�vt��9�o9u��D�+D�A޷C�Z��y�td7�3Ӏ�./�yMu��Nɰ��E��r�����w�mUP+s�&c��	~����vS�i�zt���I3��/��m���&,��:n�ǔ�9>GF�BG�m�_	�"�͹h������Q'���2h�+�`�YҨec�ў���7�WT��{Î�AĢ-�.�\QO2����a��7���P�>�ط�����N�{6ڃ�R�@�����hJs2��R��z�|]���=��$f���置k�1+��"�V�gF�؝E���VC'9���t��OAE?5�fA"N�@�>u���z�T'f(}_N����H:M��-�D�D�|��˟��[��Lh:�3^�S��.2o�B^H&��Ȥ�d�dԢ>�����^�}�����,
E�M�S�]d.��)�>	j�Zb�|�͹���rS.1����xN5�i� g��/��o�l��������N������1}�f�J�Q��D��7�(�i(t���:��x9��sq
��i��R��;f�gE
F�J��,�W3�9���+��H?�7�__���{��ĵ��Pb��H��o�h�Y;i}�@�,�a������|�����MZ�+��Δ��b��z�K�H��f|>[ZA� �����^�V��4"{2pE�<�u���e�ƴ��'�凢\jp0�;E�|��o��琣��i�P��z+�]sp���&vtHl_����V3��3#�	'j�>|�C~�emͷ�F+����_!���y	�.�O��i�Ɗ�o�ڥ�oo��-&`��^�[��x���� {����7�%�ɪ�э.ⷬ�+t�������ꗬ�ɭ�Ha5Ż3�'�R�G0u
!�s�C�(�C6=��٤N�\������Q�^�`�A<u�
?�[����S7:"���[��_O�g��G������[U�Ñ�w_���%��"�֡��H����o.~����9f�)���&��~��t�O��aq�~��u�K�e����BJת� r����=p� �P�Rh��:}E
����~�H>Q ̦�j�b�#v�G�
q���q����q'�_Y��vHlގ��rx�_�Ir7.U`n'M��y2�e��y��z�-%���O/2��x�ޖ[�\s����EJ1����n�n���Xv9Q�#����]�b�VA�����8Se�x���}��?��|9�d��o����tq����静c�N{#�.�+�}��Q�5c'�];5�!t��&I��S��4Y��)gQ��,E��o�`dQk(�i�şڶȺ�'vg׸q��/�e�]@��K�gEP�1�԰���N,�9��k%@@�:��瞌�i���=��&���oA��u*��{>J�'��	fm8�
���W��Dz��^J]ء��y�����f|b�3��fxwP��G�Ӿ���o�O��:�������Y/��E�Je��(�r0�
�ɭ �Z�72����e5WW*
�m��o`⩸O
�J}�g�"|��]����[���%Za�zJ�Q�B��lSf|�>��6X����veV���7,Hz=O�L����&�����[���&?2�f70G��WJ�����Z^n.`�c�@�����������س&o�r�1����ʃ]������aV��~�ovCB���3M��`��(F��,"aѬ�T<�؄BZm�W�ԭ�y4�?I��~���-5�JĲ`�ez+��v�=l�#���3�	�Lʚ h3+1\�f��K0��<��b�h���ML�+�ޔ�֪��x�H�2�]��p�x�"��H�O^�z|�?L��#���j��ۄ6-X���>��m�������.� !����Vʙ���a7��)��?f���%h�B���)!�5�oB������z�{��$�U��ʝ�c$=7����+`�xUn&!;�uJ���᝽��U��1r�i�nɚ��^bU�G���g=����q��n⫟��ܮŞ��u;�R��T������z�og���D��֎�7y�s��l|˛L����߂x�w��N���+ Ϙkf��M��1�&"Q������!P��d��]oKh����$�������B��:b�D�����y��y�N_q�W�Uor��e���;I�����)l����������=V'r�z���G�"-��9�H�����w���!�)*{���P�V�Ŕ���z�"3�v8��}.'@�zixMrJ��Q���40� ]��(}U�[��R�ٲ���{�:_�=�]�w5��/�F28�u!iL��1r��e?t��2X�<���.[Vr"#e��p$�$2wf���갛'���؄Bų۴e��-�$~ˇ莨��Q&�-�F:@g:<��̛-*G���Ӑ�J�N�p_ݳn��Q�mRs^RP�p���X4
�0_0?<�u-�0�_�����z�3�>���vb���u�,s���c�̳gk�jR#[ZR�v�>�duaM�ޕ	����4�d��j=d�c��	]B|��k�-�������b}�ܲ_������}D���%�1�ک���]���C"�K�70����j�)<���Z��.e5H��8Qz/��1R����X\T�k�0r���6��	��Z�ȥn`�		'	��+Q���}r+�j%�A�r�a��g�vx��~]#�J�N�ݤ~; ʲT���|���|�ţv��۹]p͇|�ћ���FS�u��&��cc������*��5:���DW�@��<�V�â�����0���å+��(p�4�N=��b
Rnq��?(��Jv���C�glZg�/�Ëi~V�Bh�` �k�����|_Y�U�S��N���W=Z�{m(�Zr�:�0
�!c�����չT#��>�>�C�{ �_�n�6�-��G�?�
��f���z?�3>����V	�<m#Tԁ�`oIM�9=R���Pw�9�l;u��
������S�-�3�jA˚[��O!� ��ȁrCB�^���`w����~�N�)'�M߷>W~7%3,�sj���RL�b�A��Ft�	E�C|mF��{oI��i�7ڔ��3B_�À��ʸ�Xd����"�"l�����r���HOo�V�DY�}w�#����6�6�N�7ͩ&}-���V1�V��q�Ɵ�֬�(j�����Q���8������si�xl\�4���0=^�U|q{)Vx��3����x����{���%^�]�Z��ݩ�����,I��ǟI�=�UӶǫ0�R]ƽA�'�.|�.�I���=NL5t�~U:c��&	9�3�u��=�>E�QԠ�ssVKP�{X`�uP骽|,F�o� =H��&���>�|P�\����c��pX�p˪.y�s�z��8�)G̻���>4�v΃Y���'�RL<��'q���"ԙش�������m����S;?I�&QR�u9����������fďm-ы�"��B�p�4����[0���w�{M1�񟖖8�O��<FHX����M_����(��P�YBPc�[�a/�1��}k=���\�$��jL���}Udn$����W}Q2��9h
�g���+�#�C�u�N�7:��S��O���hL��2P�9��!�pZ�B�]���)�5yXܓ��bG����6u=�G��Ҷ��5O!�#��H�M�R�J�$�T��r:7z�\�����j�l�T�pu�1�ſ��%�M�wS�e�FBW��+jC1��%���,�u6��Y��7�g�jGf1X�/�C���
^x���6ǎ(/�t�x�]�Č�ҏR� �%>K\VV��K2�ə�J�gg:J�
V("1�i�Z}N3��&DE�)�����4���G�c�<��p�O���,X0�H@̓�����C����	��Tƌ�j��D��	E���
%���b�����J*w�w�}�{����ΔK�z�nxt�o��D�C�"l�#ޭ��3#��v!V�l�s�����!:^�� v7λ�,'?�o��jO>��[|�	�:7ѕ?�M�O	���\�?���J+��ڝ��w�\�}���1Pc9�i���PN��&N��M!�y������pm,���{�ԋ��=?5�(�G��z_�jԿ��FU2����Z� ���C@�;j{}�O�PA��%�l,/�z������+���ܼ�K������x�-	�:��l�4$�bS��G�#N�N�UБ�����B�t4�u��k&ˆ_�TV��8���?-v�}<�2xN��蔧���x����<�ȡq2����b������x/�� �<�,W?�g��/*/�5��m*]�V�J��)A$�{1S��$�
�F��~c>�y-��_2��+M�0��4�'.\>����ŷ��	��6�"\u�nO}n�F�$�}~iݵ!�_�U�t���_�!������g+��g���{(w'���a��.ox?{�O!�K��I���히����h���'W�MYт�p����F�O�#��ʋh���-U��I����RjmSsX�:�Ze����	;X�F�E�4���;��%�H��
�����ғ<�zw�Vi{gG�� $}���}�]_Y���6pc�����s�-M`9�Ek@`=����-�H�P�	*H�f�b*�XT�Z�$�@'��Be�Oh�^ɬ��R
O���H�.6g��#п$�~~)���� @��+j/����M��`��:��>�&�à��gNu�l�ͺ]�p#������ݸ�65N�����1!>?Ʃ_��z���3r�Z	fX�� ����;�y)� ;���E��T�!��Z��q������9�ѥ�[Gք^�'H���N
b��X6L^Cx�L��(�dc���`�,C�Y�M�&##p�2�"�u�"js�q�RuGb��j��eW��C�~n&1�Ԟ1+13��s���pb��oؐՌ�^
��_���X�̂�)J�#��Y|�9�P�"��7�/���	h���:�,��ן_S}�P/�炄70�������3E�?y�|Fm��2�i���Z�\<Tyj=����aA�H4HBY��HzL@>j�8[)�'�ɱ�#��P�S�ÕF��y��:B�2������)�5�����`ɞ�on�F�f� �d�N߭���BY�{/�b�m�.lE�R�:��}3 �J2⡜�R{]�ȑM/*WJWm*[��(���z����$K�q!��}������kv��7�v=my���n>/��z�[�@!��-��U��_8�qo���i�p2�$���%�N�����pĄ�L�^��U���m�d�Ѕ^�@B^��d�vC�����=6q� �HO�ЧGޥ��:� {�Ƽ-�ob�����%	��ڛ�Jٻ��'߄9�/��>/��>;?����M�fA�9���� 	���O��!��&	6�J�1�'c���h���T�^��"<e�6���������.����ڲ�S��0���{R�: ^܎ܻG�+W��'3�ŷ *��A]��<���^.B{�)A��g�Ō9U��7'v(�r���h�^5ϕ�W\��=ºUH�J�v|�=�9�&r�������Kwt�{�H�����E�&�fG��K���NK_:�N(}� �����x�V���p�ۚձQ �K� /�e�5��V�q�՜�q���b����H��RK�����O�n����Wsyֱ�<bp�R��O��P�eh*���-^cjxQ���J�	M���"||��� g?�F���%���(Zg�_`a|N&��� ��Y�]Ð�m��7aE����|�y ��G��+1T���[@������r�z4t����h�P��u�`x�8y*��]�k��b	����ہ������z����E5��RJG���S�n}3�<e�&�_o�3�M�n9i�-�!�<R:��\�'&T���I3ۢz�f0�d}�	h�;�fPh�"�#�P��(������3�2q�Hd,��6[���P�����m_ƖBvۮ�Yv��{�qМ�X����*�v�CBlw����9U���.�#Cn詹�:Jz���B޺��4[�[�@����J��:k��EJN����&O��1�Q��q�!�I�*��\�F�9������W'�5n={դ����E
U�'�Uv:2Q�&��σ�듊��E4���p��!�Y.��`St�v�����_4�0F��fx��׻�)J���~��D]�_-?W�o_Y4"�G��[�>2��_��y���}_��q�Y�&�sh�QRh� �"Z+�^�9<}�8ŋ�3c�����`�g��6K��O7mw��RyC�+����+�8�T��j��q�|�՗TVs���Ek<�������[d�ر�Iӡ��ޤ�4n$�С�
G�J�EPS@9����;��zXn����<��ܰ���Ќzɝ�1��5�`�������L��6F��X��Z�~��t\~w�3u@]��(��7���H0�P&}��:Jh��+�o�w����:8�D����#��W]#K���y�o��(�JI���}�ȫ�j�B�+��pw �r/�P�$4�呎���_�s���8p�,�&F�*P�E!C"}��
�ja��V�G���\�6C�@���V|E�d��@ق�J��_�*.����s�"m���@����M���2S]e�8x���K�Q��$��qz��(�H,�Q�������
R3xZ�Ogj�R�]�������p�}�Tbo�U ��_�v��Q=���	-�8ol��Z q���ȿd�{7�S�<��u��?;f�����_	�c�P���7�L���@�t ��4|!�\��L[)9�����+�h=��{ӌ�M!fv�:�r)�ڧ�C�:|I��3g�oB#;!�%�f|'( ��õW�l�L(��5��޴PPPH��G��fZ��}�g���Fʨ7��a+�?zDG'�@,Xj��m��g�z2���um�����K PEF�OW�3K�\�=sU�R.�lx�=��:�:|Yǹ�M�����p-s�e��L���n���<���5��csu��_� �����]{����}k-�h������N��}baH���iT�a\������m�T��E/��E@^�#I��W��^����aW.}��+���:�$%�.[#�^�љ#�ٵ��o�-���ّ��) ��-����٨aJ-!��+u�]8٭O���sRr��E� 1�al�	�@g��S���M��R˹��"�#_�{X%]I��h�����"R�	������H�۳�O���	�~պ)F�65>�dU�h%�a(s`K�4Y#ѡ�T~z֟���3;�����Rv���Z%0"w�,)�{�3g�h��E=���g"����!�7��!Pv��H�<k�l4�s8 �0�B��~�U�zzz'B�����.�u���9��K�%&׎P���9��kx{d��&ee�Ҧ�E,>�\`\fz��e�x#�P���Y�C�!),�5,���'6u*Hߖʉ�9(���&"	E�}F��x��/5v������ҹ{�<���� Ŧ��*$,��0eU�U��������%��o_���������ڻ���c4ɬ���Y� !���w5�D*�`Ń�Y˅N��N���*���Gk𑹢")D瞴��#�NNT9��Zj�4�VR�����c`[��!��� 
����P+��Fj�7���,�#5(��%d��c�V��f�<��ȫ{!wsO����G��![���X��ӯk�#0!����7��_Ŭ��84��Q�>r;�V!u��ތM�r�\]�S�7� G��e�m�\�=~��l3Xr�9��8��/-���~X�tU��ƾڙ�\b6�>�S��	��4��Iʹ�))��N���q�������&ؘ�U7'D/C�C�
��h�ܔ��	���;�g���I�T��������������kYk��MR��(�Kf��`��Q��g��y�:�m���D;
@$��B�o��[������^}+:"�;F+�Z�O-�$U(�i1�`*�W	ޤ�(���ʼ��ݜ�8�Y�7����+a	�{BڃW{�g�A�U��a�˥�Xi��JV@����u�h``��
@�)޴�O]]]���	�{0}�#q���yJw�¿y:�rx7���~��/�4r6^]�f-@�d8.��8�e�p���N��L����F�Q������|�t��M���n�"a��U�OFC��2G��5&� OW�E�>2KU���ѓv���k1��ɔ�[�^]�L��&�����2sҶ_^ˇ�Z�ä�D2����D��[5������߳���H�nM�6�1<}��яxA�s߭삥l��������9Ě�$�=bDfx�g��=�.���@�6�h��k3w[��	>��P�l�����Ț ®�Y�q%��r.��}�G������9}Z����dL�/犧�f)�B�k�&������Uu�QR�9'��k�N>(b�ni�����c�V�U瑶`��E��1��Г"��c���Zt��>[۸C�Ѹ8Ѡ�%��NY�ϕ��\�� ���G(��ܬ+�
�8����o!�l"�כ���Q�?%.\�s%���gĐ>^�t�z8�~>ﱮ�٤��3ܮM|�-{�>G�O�c���Pl�����M'�U�g�WbƂ0�QSQ"b�b�f�0WH\*����.�L7AY�o2u�c��u����'-���
����JA�V��<�H�~�Q`m��X!Dl(vZL8Ś�����g�
+��<�豅w�yK˽~g�L��*W��/�Ap���D��e�[^������Sm1��]uj��*u�7�\h+ŋw6�(����*$L�oE]LI��m�Q_;��4	�u�J�00ݤ��x�<h^�c�J�{��Ԑ�����y��n<�jp�_����1�^�5���i��Cc?���B�V@�Vf5�tm�ITPE���b��}cK�u��d()�k y��b>�n�W,^x�1���o���@WDu���sW\���!�@�υF�	�1�����(�X����ԃ�7��(�o^|~�K"�K vt^]߅ф��̋mD�UeX@Dg>���j�Ȗ&��s�؉���|8Y&��5�%��=���>`����h�0��,z|j�����z$8^��LDt׎J�q7&��y&�Gndk_�����hLܛ;��|m�;�NOpԬP;���m��,���
[��m�}��
U���=h���c�@MG&d��P�_G�ه[W;u�B B:|�=����H��j�]jG/D�4�6�~��L'b�&0\�Zl����&�T��t|�פ��w滰[�ߌ,���Ś��~Uh�$K{Thq��B��R|
C���.��h�+P[����sQ�#>���~�e�t$���;e��vV
q�u��[�s�Ƴ:E\�(�����)��_^��:E�/yeX��I��(��Mtڸ6�w������ń|Jʤ��K1o#��^�_Q�����]I�||sJ�����/1�׮(��q^�1մE��OO���3y���[u�&&�-;}��y��tK�`���M���G��4Z+�z���>��ܳ�Y�p]��.�YBF�'�k7a{t=�'Nk:����]X1V������W��ui��|bi
?��y�u฽�&}մ�4f\wR�7��x��3+�3	��ң馽�LY�W+A^?d/E�`�h?(t;�r5`��"Y�'�t�H�y�:���;�ʆ59\�w�S>�ں���D�E�'�����9�3Sf#Ϩp��8�\�N�
�ՈY�3��2���TS�AeuP�=�'����W�zcST~Kʟz�j��b9Qr��	؁�c�m��H$�f���#cHB�S��]zRC���͙�-��dP8��Y�Ǳ?B�,-ŌU��M߭�xS��R?�t�����9<�9�d�N��b� 4�./t5���E���>©߶3:���!�����'%4����?܏��a.�����nЎ����k�ҭ�]��JY���wS����+�� p�z��(~�x~wn��8�z�'9��Nn!@=�KT����$Z��6Lc�o�
;H���qQ
�� �ţ�h��1[mrX��s����}��N/$w� ����:���('�@:"�`���f}�|5h�K���B���u;�U���(�B2�zi�$�{@ā�{S���}���jF��)[�]�n�"z�$WĖ׻�����5���������]2�-/�.lj�T�ʜw�̶M�� ���]a�S)�c��/�)��B!�h
mX���_�8�Ӗ�H�hn[�|\��v��j�_�89�L���64YJ�?v��g��{1�����I7G����H�]���YP]M��J+)��	��Ĭ��*��ϒ&�%��������A5=+d�}葮�J��>�`�=B�c���f�$��eY�{_��j���X!��{��7�v��8��{�{액	��@[>�{35�1���lSh0 �H}�<v�[3�r��{Otl��aOSWU��Q{��h��ZP�Xˑ���C�������B��_*s�x�z�_av���a,��^%4�sN��;���7���5 3�.ĬG�t_�c�w�c&k�x
������
�£��;έ��(�Su< ���!���F!�����̛���'a��F1��Ȉ#���Ο��=n%�9S�3e9V�����t6ֽ)��}�D��5� �'Ħ��)@ה�	��P섹�������^/��Ƥu����|���k��{�r/�|79]�V��d�A-�o�`����x����+����ӫ�4ͽ���k��Dp�sV_AV_��l�z�@�!�{�����b4�[F%�E��u?�$y���	R�R_]����o����Qτ��Cz}�T:��U(�k�5�e_�
J���[u�l��B��$eY�gu�ǜ��Ս��	��\팩�<0\�������8"E�������#��\n[(H&��T�0�B̥[�"�î�n����֍�K�'a�q��� }���e\ۻW������e�ok����߯�9釗�>0#�������I�\�p-��{t�� |�g���F��������)k[�&�/��������Su'�
���A�O1~�"g��j���}��[8W���d�n�U\�I���7�x"�H�9ku�Q�VH�*����׃�]���p�֠�_CS���h&��6�ȟx���k	c
���0��Y	`�a�L��I!\�N��_~#��0����~A��M�H� ��f� ����W�����Biqoq�BѲ��[qwww/�ŋ/���N���aqw׻��?�>��n��$�L����t�s�b2Q�#�X��Qx��k����=y41�%2B����J4�'�C�Q���*�}I��A�LU�0TA-����w��-x(">�ST|Z;�%�u�H+~|�H�V?�R�Xѐ�	����5�P�5��2,JĆ7��:A��1�'�凈[���e� d���F�t.����6�Sc�D����Bwc�@G)��B��
�}����=iKW"�,	��X�q����5�i
���J��Ҡ�Q�,"d�?B?��B�v���~�KA��0#���i�fDb��!LC�v�r)Ɇ����V|�Q�A�c!DB�Iǟ�����I��
���OB��7Y��
b�ؒY��V���-`H2�c"L]j�Яj��$��bd<X�Syl�K3[�C���'md�?�e�u�ewCׂ�9��hN�vfO�mi�)y[ٹ��!����H�j\����&����[�9�p`��c�� �� ��k�����D�C�x�K����T-���4����!>ABCl&Ͱa"@m���5{E<��H���6H�� 2��͝%�Z9�q���X�|��B�5�8]VӗcSF�j|�5(#T��L-;�b	�b0�I[�h��z�.i�c�jw��9���I�Ľ=z�`�E��T�k�����C����3��W�����g�������CA����O�k�l^�.��`�>Wr���`p��y�w�fF(��_ОWH�N�ډ��]�bȅ���G;YD����m����8���V�:Qß��i�-��*�/"�P���@��y����.4&�QwOnI��+y˱�_'=����h�.�K+��>�]�+�$e�(���6�e��ʆM��EЅ��6����D�S'�"�'/�~�^f�	�h�iȤ]�����b����A_��U�H�%��r�׸T���q>�p�=�
���P/��Cg� 1�4�M�
�g0�߿����6�ӿ ��N�{+y�V�4P�R�<�P��5yh����E ���҈z�|1�x������J�{&0�{!��N/��<+S��ID''��t	���-�{�wa�1��յN�(_�C9��!������խ�B�cG/��C"�.">h�X���=a�X�:��?a�D5���&�ˈ�7�{uB�)���b-e�A�.��m`r1�8��f�P�Uw�B7�5��n���M�CY%������2�4r� |�"r�:B ��Vɳ��݃���~�/��9�[�O�d�*��M܌=3�m��ỏ��Ι��aF)�ԫ+���q4�k�b���+N��n��W�ϼ63O�i��Wŭ�Q��M�4;9�
rs:U��jэ<� �_E�3��}��H�ݭ��ن<kk�6A�����r2��D��?I�a��K<�r��2Hl�J]��ʅ����Q-{Bìy��f�*::��6�b�J�G9�b�����؀��U)��:��|�<O�sX�h���ښA� �i��B�6ӵV�v�:���R�D���>�a�:����
u׸&���>�Φ!0��r�� �`�l��`��0˯������2�2���ھ�">'����^]�$�C��>%B�F�Ђ��YxH�Ƽ�b^�[᱋�C�������������:]��q}OB�:00��n���<7�����ׇ�5 Y���9�;/A,��ֶ�B��g�^�Q��`�ػ eZ�����-��e�:�_�[D>g�_�"6
V$r�zy��T�W�R��t�ڼ�HKX\� �R�`˽���8Q�7�/���T���BF0:��{�>I�9�e�%b�K��
]�����ڸ�&)p��D���b����]_�-t����D�x`�;��͢���F�ǚI ׵m} &K�[��z����]��
�Zr����#��J]ս+B�׈���]�_�J&��#�m���n�㥥&�_Z<E)ᇆ�kƼ̩�wJ��(���P�	�E#J�]�l�;��i�@K8�u2����'p8��u}s]`�$ը���p�{j�>�_����T�A�TK���fo+s�'�B�=�E	�;D�Q���9Y"ϒ/�C/1�<�9ĘO��5�}9T�-L�<�u���yg�zRI��r���\���qI(���Lq����	KښF�M�9*f��}.yD>�Y�_f��#օ|��Vq���ej�q����=��F�2i��j�B$2�����8lF��a���9~x���}�w�s�^+��_:�$���T��2�c�/2���,���Q��Ĉ�@�H�b��>>d|}g-��k��?������$���N���dK����e�t��������n�k��F}E�웏ܰ�l4j���D��%��(�ƥϚ��K��H��)rᘠu���`�vz�Kt5ʶ�*F��yDغ���~Iy�x���1�?tq�{19͆;`!$��R��E��!n],��$�}�-&}=�b�J�v��(��r���s�m�|i�wdC��m�o\�WE��l�������ߤ����x�1W��(�z���E%k�����4׋jB9��o�T|��=����#�Rڸ�F���3�txϗ'�.���?(�A���/�b����rMd~y`�da��z*��DZ/n��Lh���4c����J�I<υG���ޢ��)�#4{�S�7��V�۫�N:�k7P��Ø�s.K�v�$i���+����f~��n���m1Czz� ����1�;���w7�E�2 ����fZ��%x=o��z_VhȊ2u!:x��9�뮍��}���3Ѣ�)��ͺ/^:�M��=���5���7���������D��w��y�X������1�iI��� �qPS͆��
�x��T�sM#���$m
�ʦ�)�J�!�T=ʝ��f�9�q�ŋ�Ih��T��b[�}9� �#t��i#3Σ-l-Ʃ�R��c����e~\�9"q��qz� ;\k��D��Y\T����Rb%�W\����i��ܨ��m^~�E;��}��0��Q���Y{x�Ʒ��}�eՂ���b�,#��[L�"�"��2'b����� �M�1g��ݨe��3@��βʿ�L�h�.��ƀ�܁����U���8w��`u7Ԉ$����U�GY()�s�Us���x;���;��0�u��ڼ.QZz��z���c[z0��o���}�����L�m{`,���5��2�ո�򗢸�]�Pic��gr.\�T�����>ܰ�}�O�T��^�Uy���<ĺ��>QI{�QMI�ؖ|BVX��}��
��[P{;�ZW�ɊW�Ǐ��^�ŇT�:��uWo�m�����!x��}Q��fK�?Գ�-�D|��v,��.5ĆQ:n�&٢��h�M� ���w��E��/�w	���4$`KzקYD�d0��;��>rt0�#K���~�"�di%t��������c�A;�[��3q��p ��M�Ǘ���ː����7G߫��dzBK+�eĽE�w[vR^a�tm�LU��1J�ǩ���ma���E�p2&i"Q��u����2�����xj%����t݇ܢ�o�?�&�%pO�g��鿡LA�%b��YеwL-�)DJTG��_�~�E��i"�Ø���t�yO"g�+�A�	Q>ƃ֢e+y��9���uKB�r���
_�������~%;G��|S��V�������uЛ�z"z|�B��x�����t@>�B�rL��?���׽`"�t�E�ה���Y��)��0�D�p�ˏ��R��`j���.{>��~9�م�u3ݹX�B3+�b���� �������߇3Ø*�xw]������oM�@;�Z���1j�ob���Sb!ɨxy8�s>���������˶�v�A;ً"E�wJ3�7GϪ�	���u��j�N�0�ۢF?x=�hD�Y�+#��ޫ�� |4Y'����mL���v�Lo�7Ӓ�1v01w���\� �
z�������b�o�-W
2���J΁�Ԏō!G��=X���BRYC}�`���:�w�D�Pm ӄQ��K���'ڠ�;��I�a�a�|��0!{O���Z��ـ�h�PX�p(��kݠ��"�r>=7�s�+plZ�k���]�ݦ�����)�oUIt�

�b ������mN~����6�C��+�)����5<&�Μ�oGP6�M�6���
<۴�w���n�n8 �NZw��H$Ы��E�I�&.�:��]�<��u~�_�e:��j�5S$�!����Y��1�uwl�����>��'���4:9X�-�a��W�3Os���CW?${4A�X#��A���z���ח�{��������T���/Ws�Zþ���BA��@���U�+ܖ�t��oZ�/�I��5����=���h�k��|�ٟ��q�����,��!M��Ӑd�-�~&֓`�vx�U ������l�S~鳍� ����nu��z�Dzpo����w6k�{3�9b}X��˼�-�^H�����C��+}�&�S�'����A��������ϣ�:<��W�s*L�'d�S���m ���Bk�������;uV|^Ŕ�sv9����7��n��4$��F�i��z	$�:b[@"�p�kt��8�7�ji��l���)R�1�x{ �>>��7ݠ��}�c�`��8z�>��ju�^?�V��T⭅aѧ�ep(�߾�<f�����dԫ6e8(���v�Sx������\�Kw��@F���3Te��i��(QuW�oxL�v	;��o��b�.*���6^8j;�yY���`k��	�Qv�W���(E�oSk��C�y{��l?�ɋ�P�����T��Q�cIVgҭ�����ɩ�������=�X�q��P�O]�I�¡�	��
"f�K�[K9��c�ン�&<D'��?B�=�vl�����)6a�}�h6�|��ǯ'���-,�Us����P2�yG,T�>�U�������+|QKC)�ݕ�����F�Gӆ����̖�W���R�-çu��um�i�'�꾯{�@��ͶU�h[���+��n�AG�;���������$/�)\��T�_A���Q3ѷ><LѥP����r~>��Ir/��ٳ���<zx%���<���r�ɾٚ�q���3�C$y����	�F@ۏv������?��mBy���Q��������9
Y�V6��I���>Gi[�B��a��Ó�*������L]x�
�*Ǔ�{�H�3�N+d��ubX�D��s,���ۢ�%�y�h�2fUC���i�A!.��pz_4�Vb�#������ok����
�8�����b�i�5�>_�szU����G\%?��cK�SV�)�
'd0d����r�#V�ǉ����|^
M�X��_�!&�R��4R�w���.�����>Z�c_鷺i#�@�)4�L����M��!]V�z�b��h3�)3�����v3{CC�vF��V;F=W����A/d�T����罎�4�K�Z2߾�?�y��(��0[���E��ﵙ	��nW�70NR0�W�_��b� �d.3\(�#,�h`������X�"e|�k[2��y��e���Z����kPAI�F�CӀ���)q��՗2I���O��yQ�3j{�ƌ(���%��.E��b�$8���T���X�S�0H�'V��!��2�$<�7y��\��b�u [����E9�P��6Z���c�.�DЏl�>��ў֊{�L��j��ͫ�}y%_X�����7���G� ��a|T�0��,b䜞�z���X�g?N�^њ��D��Z��E�.�Q����a����7[80�^�3m���Q��h�$	t������e9�ǵK�`�A���=�͂���������7���RX��f%p/�i3_�q"?�B���Ma4*�wš���g!�����/Z ��f��|�m�
O���8=�[�W:���]��}S��##gB(�;��[u�(�;�1M�Uy�L���y����+4E��	��en��>8������)P���9�~,���/y�b}<�粶L�e�M�-M��7v������������ˀ+�������T��Ə��n�~w�Q�p��S��T���e���!��k~�˧k��b�mJ"ڑ��;t���N�6�}n�1�;�F��핳�z|f1�����r��v��v��U�1��nN��;�;I���g	Ft��K>�4�wՏ��q��P9�-}oé�!-Zш��qB�y� +�7z�J� ����yMpJ���K.�P�U��~M:+��8.T��E[P��P�y� �\5d1wI�}���%�,���I+��g���㈖�j��Z����Ȥ��7_Yf�Wٗ��f�����o/51�\�����?/s����S�xV<
��J�ӯ���
��%MM�N��oi��h���@���C����&��v~B�>�d�]��J�<KI:���0�bZ�w��	E�9��� ^'�-ɺ�9����������f4�$3Z�_�?I����!�mh��=�c�S����,B����R4X��������m�e�����x��%?Ǟ۷��m�)�����8��?��+��Pes�fV��쐑�JE��"	h�*�~�卶-E�u��Qc�=�%rU���#$��s��uY����~�g�����i���o��]8lπ���KUi=��8\�����еy?f�2ቑ-z�H�bתJo�}{����lzTl.O3Y�Q�>�%��b4�v�8c)B-!�ԌaqKa>�� �ߺ'�
�5m�?���t�Kk*��{�?'g�0��G���O����)_����Q��LN�uz($\��b��]X;����%��:-UG3Kŕ�WdB7��w�O�	��
sF�S3�=oҫ�����5v���t�(T4�M�\gfs[5�Igm��9��a.nm;���*�>j++'�R?e��~��z��OM0�jV�ej��Z�I���O���J��x;w$�؊wW`IbQ���,���D2�S�.�h)�٢����b�H��:ߔ�u�F�ֻ2�mz�۾�q�d�LR̸�QZF��K�ZZ��u�6	�K�MӪN�^�+��A���ޏTIV� b��@��C�t���h:��@ö�����ʓ��@`*��V�:���Hp����!���D��Ŕ�6ɛY�cϼ�x�Y���;*9���2G��_��hq�Y.�ܟ�Hv8<�_��^v��"���Z�e�dOtV�mE�����oR��)�+��x�'��D�-���%K��z��Ֆ��$���ѾfW�$�>��(�*R�RI:���|r��@�ۘ�~��8�"�(Y�l���Yi�C������]�f�ȝ��5Y]ֈD3��w^�!�K&�Q��K��A�Zdr�
���"
��ӎ�;��縥����%T�.6�dt��ґ`5^��H~��f�C���\]��p�2P�;i��e	J�<uZ�5��+3���I�\
�a��QEd$e7���t���D�7��K��|Sz���;�vQR��Y4S(cy%Pt�(}b��
?j�텶�т��^ꔙ֜��D`�j��퉥���,�&N&��F���/4|����S�����Q$�����}��/�q�$14)c�$a��*0'����擒��i�߭�p܊G�߅a�=J9�+b�.�x>Oճi@�CWQ�7���%�a�L�6����{��ͮ���d|��Z����~�N>��}��a�?6��D� ���w��}��dGΫQh�g�(7,�	����f1Kb��y��D_发�SQy7p8��M��J�͸���l�����1�1�&Nܿ�g~\�n #A�R ��̭�U��>
�Xh��l�g�ÃK�W]�_�	=�;�G<�����O���'����b�I��&��$���g	b��XB~ۡs� �Cd�M�eA �E$��/�^&�r�U�&�))	�;�����#��1����o�@�H��Y�{�@��d�)<k�R���_����ن�T���x����~t_5(�'��ըz[��� ����Nֵ:���u~��O=\��n83Q9�e.�ަ5g��ɰ�0γώ�緹	��9ߊ[�pTL�b�Ik�����뭴�N�r�I����毄��A��¨�Bbqҵ������H.��'ǥ�*>w�s VN*'&(��ŵ]q�*�FðE]�=�@s?�Qq{�+��e�;(�L�*���Ez)Ӕh�n�GSn��9�?�l��=u�2k�k)W4a$�;���+���ao�'sr�6�'�������	�[2,T��_�1]}�u�9d���� p1��Ͼ�-�&���w<�I.�w泪�8]y����@�Q�핣˵�#m]ێ�� *f����.#R�z"��z�~#)]s���\��Vi��1�V��_�~϶��;⣓�#�2�����
�����	�^������!scz �%����r��z�!�F��|=�[��yz"��
�["����8*��
�S':�^���\y��~�aM�T���+�;l���:�������%�S ��<B~{���`���Մl1�a�*t����#��1�@UZ�8���Q�K��zimWI��L�S 8���u�1�.��Ngѭ�=o��]D��5�hSz2��[�4�s�{�ٞ⩈'&�;ȗ��h�����������GB����i��؎�s\)fk۱�1�����+�KX�}8�w�y�īw���/��ix��i�T|����fT��J�eR�x5���JA2i����>��`�-8�Y��ĭ�Β�h�F�͍�ƗAA&���VRw�B���g�V�?d�;�\Ќ�8`�DE�n�|d�jZ��=.���-��В9����'���Ysx/9�y��3�+u�gx���h�;��M��kE��'��Պٿlʽh�P+�b���"&el{����vz������=J������<�6Ф�~q��\zr!�"F/	�z�Qf_����C�	1촢Y��t��9�s+Q�<�<�B��_�+�^-_�W<ſn��*�<.��t;���f�`�)vH#7�s+�6O�V_:��k<����rU�3�GYn$̝!6�\|�]�\��GӍꖘ^µD0����Io:d��=��p=ڤU-�,��
�d���r��j�uz>��?���x���3y̡̬1���B��� xӧZ$�{��wqW{�{�}�o��_��8=�k7Ix��9[�&����R�V��J[�Ye�F2Z������!��P�&"�J�UE/�,	H#�L'���*��a-~�UG���?����-Ф���B[�r�}*�^�����aÛ�
���m�uN��܅���lyt�ܦ�ӻ����"���<JA���ҟ�3�=�G��p��I{z�Se!�'�"n�zL��v��4F��<��|�k���c�'�z�'���S�pÓ"���#~��x���C��Iŧ�7��Eg�fb�cj�n~�C@R�t�Ju��E\�^۷#~��Մ~:r�(l/ɜei���	�"��:��w!� 
��#�>�YPQ�>�y/� 6�/���J�KJ�e8�����3�$��B�wE#�d�����X�H�9쓤�W�ǲH[�Gp�pI> i�r����BVS]�i��yLB�&��ʮ�}���
ǚj|<{�����w�P9[	��F����D�g�ZhVQ�]��6Q��f>p'�I����|q�
�U�gά���Q��&Ӡx��"M%�)���4b|~#�a����KKLz��&�o+��\s�'�ZN�q�³ʡ��%2����+�g���=-Շ!Y54.<�JG�4��vzB�����j �
sHGω�l���8�[>_�J�������%c�4狳#ձ�������/�����F��d���7a"z=|I���ɼ�� �&I����9"O�E���fC>�h�1�-���s���4��<4b���<�L �"X��:^>QC@r0�#���Y+�~�LPfA#g��]C>[�×`�_&���,=�_�ꐞ:��}��X���m9XC�&��q�*���{�pD�ô�O���T��ι�V�:�9Q7'4>�$3�T����
%�ٌ�~�.�l��$vSԷM�e��ܳl�8�UC�"W8�t9�����4�ȯ�j�@k�#YD��nj�Q��2ʬ�@�R[%$�����E�_��ݎb;���L�bV�N�с�>7��s��aܯ��ߋ�A
�:�����?#���e���|�;Q5�'����4�{e,[GJ]5�p�\~�p�1�P{�)A_��E�φ�!{�Y�ȧC�*���XS�oIDd�x�J�g��t{v*B$*ltr�˿gd��f�a���R��S�5�I��u�'�%�Z�=���U���`��,p>Cp6�a�|U
*b��>ѹ����g��V�,_v���*/6|�l�׋��B�;0|Z"�2�ّua�tbU_*(g �J4�)K�v��9O��%�aV���m!�*t��N����ɱ���K�l�y��j�.Ǣtb�4^��R��e/鬪ŊO���:���j�v�Nk����]V�)�2�Y?p/`2볬�s��������c�g��oe��'�P<�Vx	a�m�V0s�ʇ�~:8�P��e[!���� /���\�%Z�kU$IO�CC<���5��(�ZC��˘A�GK1��z"���yH�9$5�r}�<l���{�?��0�M#@ՊV��Hia��0��$P� �b��Z��E�A+%���r��i\�7�|�s'8pȋ�A"w�b ��K�5�`p�[�k��W>���%Wu�(�С7U���I��l�%	0�������[ߧÁ$̝�ja}�m;�9(��@�4ӂ����=�_�B$������kQ�Y�e��E����M�9O�!�U�F�wD*�o�!�%���X��J�/MfĜ�HxS�=����T�QI�L�:��N�U26ӄ�r�D!�z�ؿ!nP/�7BQ ��Mͣ#��I���кwm�<<��U��`���I1y���m37?��&A���oૻ�V�����7�Μ�HA��� 
"ReP)�D�6����|��-�i��Um�$��|��ql��L2n�?��޲��.p�9H����[R����ԷJ�(b�tL�tD�R|;�=��QlX:Qe�g��^���C�����I�V���L�o�8��n����L�cA�-�`�fAK Uq��Uh�i�~�PI���k���ߪ V
�g.9��br�����[x�\��T����+d���6�9�f�M��`C��{�I��5�[�1�l0����(Y�$�� �[�\=�r�~��v"��xq5��Ⱦa���@� I�#�wK�D�y��P�DA�pA�Cء�Ǥ$�o�W�o�&��������K�W4�`('���«������
7�~��-)��������lEE�J���/�9i�N���II9J��Q(�F���"�9J6�oj�I�ʥ�~�
�b�G��J���v(��X} !jC���r� "}t �I8�<p�'����ua��=�F�CL
��O��J�f�uST\�Ҕ:��PHS8D���q����5��?�E�!ʙ����h���~�_B9�>@�����
�MNo�-�b���?L�@���Ax�
�u`K���d���A�0B����Q������8a���Bd������j������+��Tb�H �{ߜ�1ě� ��&��}�,���?6��~̡ˆ2}	��`N)�	B��}t\��s��M��nZR'SF�TiH/��O����D%�)�ӱ�e�6dҁ�:����@��Br.J �q��_��!7Q}0�5\��!(�-a��7L�<ԭ�ä>�/�ǤnZ���G >�<�Y{���� �Y��5?,JZ�*_C�x�&1��j��=�������+5_�
pѴ�y��n*<����$�^z�33ޔ���B����V@'��`0-ܩ��vL�(w�N�~�
WI�Ac�9����P�D���6BV@�����XD�37$�I������i�4M`���pe�����>����tN
D��{� |�����.��͍�n���`m��B�
W��ED'��'�P@���yz�2�2ƀ�����0y���v�`��I\LG��W��H�_���8/���(��#��B+R;����o�s�V#&�?�ג���V#��X���='ix����	~�c�m�L�܎�mz���B��tc�`��#����x=:���ٲ�c'�<�{���~�!�\.���H�+�{��^��ݓ��A�7�۬�'FJ�Ӈj������{�F�.�����Q2e¯vwnI��WT3������є�1�<[��M'� ��;(7Ǧ�t�B�.[��GW��g윀�Tңʩ�]Ym4r.�G�_�yj���z�y~[L!�r�̄1+d��c�I97���54�@�m�͓�l���j|շ|��|�����3p�b���Fda��\�E�m�_;+|F�9�o�qj�7n��O*���C�x��'=6��,�;4�/Ag	h8e|��T�d�.��~�Q����
��&~����|V�c/�1���#To�(�\	Q��J^4�z�W�Orҷ/-��3��c�[� ��4�q����v<��^5�1�U�AH{�g�ڑSVV��n�{]eu6��D2�#^�%�usQ��'��#���Se#���GK����ƈ�P�2J���a��5V�\�Lf�g(����٭Qx��b�Ƚk�9�]@�V����I��ĳ!8=�;���}��6t�׭���P�KV�=�ي�;���!-D������"���a��o���v㸼��ݏ�{00|�FN�^vU�YU�-�hq�BΜ��=��{:v���dH��i����VSu��?�-�x�E�w��}�OJME�?���IE"�g��=�Rs��s�4c�����K�q�TtyѼ'Z͏:�n���ǟ�������xp}��KDU,<梉''���KN� $�M��ښ���a�a`F�q|��}���^��[G��~ȳc�7��އ���6���.�o�s����ӿ�$�j���X�`���F�n��%ב�	儆�6t��zܳ��?�o��ħ���������WǗh�y�bb�*���.X&��>CM$*@�\|����K!�IQkG!B�B�+l��!��o���jыa��Q�s �pV�7
��z������_A55�3�R ��&��y�Q�х�a�G�I�=�,�V�͍�`]�!C����u�6#tҷK}��ϯ.a�'W�wo���l嶩��p��
a_��\B�o�Z��[C��\uCfIJ�a���������o�P������~���I8n�%uc���ip�i�ӈE�^�z����Q�~Q"�G��&���XxH��O<>튟o�u�V�c��m����2\l;����ﶅ]b?��e��C��=�4�$y��L8D&svɏ�$�y\�b��E�9 ��Zot]7J:�T���c�yI�>�_ut�R4�p������ڀ=no���p3��
���XM�ODC ��p\��"�K[ё�f���d8�4��	mI��3���3,�Z��h�ր��znM,t�|{��Z~FQ$H����D��X�yB~���9�f�8�Y�x������.aT�ƥw��p�yR�Ǻ��Ǽ��dE��k�2��r�F�i?�k��z��1�_"#N���H�~5�cY<�.�%Ňà�����àOq���o�n�;���Q��[��5�Pѯ��\ҵ�Gk4�z٭Y��F����$�j� ���������'�"�����R?����o�sA����I��<�w���4�����x[�q[�cO7o�-�[/M��§z]���b]��N�୆�Z�����B�ʺ^��W���,g����o�{^7������^mz�/�Y��|�w
QJs�N(+�*����i�{�y�~[�����D�*ʵi��Y�D�*����m@.�4�=7l�r���~��(o+s�M���a�b|a�RVشq��_�~/�������g*Z���B��\�I&���!W,w�w��Ѱc�2W����Y���@�;	C�K�����-"���|������z?��ꭓ��)ۘ�2���s�/�쀛�	��ڑ��Fà�5�T���2�&�hb����߃��t�n� �>x�'4��\���O�(-�S�pm�QD �-�J�L�\�����'+��7i����׈t�����$U�9\\Ӹ�V�,��i��?��/���BI��EO�4��?d���U�V@:ã~#(��ƨ-Nz�V0��X������Z[�����b���#�Rb���t<4"�$�C�yՋ�\�R�9[�嘵,)��i(�m@#S���5��)^OiR@{l�̯s�|{&����M`�r'S��1&m��3;�����(���-�lY^��p�Ś)?щ�Y<��bS�T0����=�R��������yEr/r���?���JBԴ��R��}�n��ʫl,8$X���Y,ɡ�r+��cf��`[��&�Pt�&ǳ�ƫw�w�Ik�K�r���5j��$�pG��0�_6�ڜ����(i����8�����' ҹ�z�7^�>�[���������#�vj��^���ر��)��Z|��
X�! ���p IaV�N�w�<:P2�������(۔>�����y-�!/{N��Hd���k��º��E%4A+�25<�����qg.ԃ#V���Տm1ufs�.L�	u� Iz4��
K6�?;�Z�C���|���|[�~�U��6�C��m�7�֞��'�C���E�(y�����뾜��|��!�Kh��'mj�9v"��b��\!׼��ǀ�T�����N�.<4���>ed.�:Ԣk>v~>�Q֨8�/3/$�c`�tϣ���,��
���d���"��Z^�f�@`sl i~M��fC�&�8�c�C����ilS��\��gxlL�_��{Rڙc���� ��)�C�ű����=��򼀻:���0��kR��q�46�in&ѵ���*�t�4*�:�ѦjC0*�A��ܮF+�+}�T�˛gXd�*JN�L�� S9� :�W�v��%^y:��K�
��8!;��`�,���>���Zu[� �����W@�pP"��0�7�X��2���n�||E�B�1�K)[Q���ȧ���rK�!�9�l��r�I.����+N���YJ��Um_pf�T��u�N���饮P��a���/�n�\��8��Y��0������[��=9; .zX��Mbo?���׻�l��^�Hs�9ģ���J���_ΜpφegL�
�x��<-��=.�1N�M�5[Ɨ�e��6־@��9�Rg���?xT������VӬ3��0H@�Ƃ$�;��ƫ-��"��0��d$��C��r��1�g[��r&Z[��k���}�`�)�>��ͅ�k�p⎋o�T$��m�u�e�h5^�/���>1i+�+<�ʧ�W;��f)�d��:���2bC�=�ֻ��@�CĽ����G"�ns��G�s���,��q��n�����s�^�"R�����~ᒨc�������V�G��4\�Ҩ_��c�kI��U}n� �_�7��]l�s�ܾ6a�q��C]r4ۣ=���3��VEE�e�%�kF�	>
�I ����-sS�W9��`�
�z`k�C^�}�r�L�2Rf�M��z��_,�k!���we��'�C��xk�0�!L�ˏ�/��W���--w&O���b�uǵ��""8���q2�$�6x|�i}n�
������yI=���.���R����*�z��u>���ʎW�V�pެ/�."�t�L�h��X�9�*w��Ba[���i��O��WXG=�q��7y��<q�J��~�a{/Q��b���rc�39��4>C��xw�y�Ų�<27^p��+�}�if�;�!i�|�����d������ ��G�"G�Q&������4�ޞ�75�Jv|��{Y��&���l�kq)��9>!�ty4-��aa� b��͛��YF5˺���*-��V����/����x�/x�ʏ3[0޿�.�Bӽ��Ʃ4�ч5K����WǺ�#������t��i#.4ϖ{/��՟t
{����|�2p�8�H4�Q/�It�f8��	�Y+�^���K�"��om�*u%f;՗��|��
�<*��l4�2�3���.��r�Y��f������QT��:2L&�X5�`"O>g;h��m��xZ#:���;�i���̋�K5_�z��y=�U����:+�pഭ�	>4����@O��0���5�E&o��a��0�Y�p*������I��������:h8緬���yFwI��G���K��|\�?�0�<.��TK��D�D�6�gK�H�H���&�����^�x|K���>��&��)���G�Ti�rD�z'�=�!,L�7y�Q�	L��h����LU~V��=1�o��x�Si�N�y�j��h���p,*���>�kw$:#Վ��E��	��(l#w�Em$^ÅZ�T����8�i����ѺKr�3$n�Z����9:��mgb۶��F�4N�6�����vҠQ۶���|o�������s����s�ٗl������E�d��'��5�J����q �ܢ`�Z"��`?�@�`�/^���=/��i2y��j��Ʃ�Ν|�:?�>�}]$#:���Ƨ�Bc<O�o�*ѿs�����q6a�ʎ5��&�T ��(�O�Ypnh�,`}'�ݗ�|c����z�5Z�tO���
Del65����kf�?���V����iڷ;@�����p�^	n1�z���_�.�����s]�f+�Y��

7�Z�y�gÆw��v�/�f���W&��߲���f����on�L+%~�F��q���{v���܁��V��7d�
9Or�����=��b҉"y	�[%ϐI.��0�.T"���3��ǵ�kq��S��D���Ӯ<[0-`18������Fr��8!R��̋��Z:����M�I��A��z �ѫ
��������۔W�Fx (��~�
��������nm�(�e�	:ʠ�ј�F�/U7jm�'m,DV�T����X��W0��Ƌ���
_U�"�e�1�|R�A���lM������H����1��pl�y;���z�4�+C�ϻn�q�����@������<�h��4��qK��'���:���[{�;;� �X���
��[�����_�r�"��,��D��w^����f�8[Z�I1�e�c؟+�V�įM�e�Q��.XF��y��n+���`�d��
��.�)��v��>�KX��|�˷[D���%�9$�h�B�ɍ�"�,�
��`ɏ	^��͞-�m ��F;thk�����`����m���A��V�P��d���x�וx�C���^mv���Q1,wP������{�&Sɚg��#v'�aC��%�A�JY��)��]lWU[�Ů��@�w�s�+kx����?��/A���PD5s��[S��n�A�`���P:P��F5|������K�*M_]'R�Q���Q�!����:�^�b����.����`�,gl�rkn� o���!�7I�O���
u�-[8=?�o�4�����NE���o~�E�>�z�i@Z���ٝ�Ƿ�Lհ�5[c|l������ �o���YK�K�c@<����V�"b4'ðS\��_�A��?dY���-,ث����7��m!�޻"�Q�s8a3Jifi�M���A���l.X��u=9I���o�?��r��}�/� *F�������w��x��_�N�O��F3?��'�U����%X���)�%,�+M�O��P֮�|%a�����!������%%?P�9�e���@�<�~�b��q?�����d�����Q�f@ ��\��ɉ[P�ʩ�3�kf}Q|���a��#�f�j�uu,t���b��O��K)� I���֙ыx�f`*��m`�q��=��aX�˳
����H���`�Eew������+sP�MW���7j_ʗ\%.BuZ��s6������u2���G��%
���߷�ѬIDv�Ȟn(6>�U�< ����B%����Lr ����w���4��E�W�Ĩ�t��,Ѷ��iѣ&.�q��&#=�0b|5d�C���v�6��M��!��d=���4RH*\}>Q��U�3"As��2��/(��y$5�����g�2��ն>5��M���_]�����|���N�2�Ot~D'��ڮ}�<=�{��g��\�
�G&�1�`_'��J�ZW�阹N�xF���	�[Vc{�ً���h�r�cv�n;���L-5�~GrĖR/&�����:�t��X��wqC�F����x���/����~|�Uq�!&�7\��$R!#2Y(�F��lV����}Lkj�����9���7Ԟ�:�D��ǳ1��J8Ǘf�������#Mڅ��R��y����=�0��P�!�p���JZn~�$����9�J�Q��������H�k5�;`%
uOxNT��ɔV^9��͑���������Z�q��pޞ���.{oO�Oݒ�~9:/<Ȼ�e�!��:�����p�y��й��Bmm�;�IB��\8�wa��x�����z��#8ӆ��*�Ŏʊ�Q�pfS�V���k���*��4c���?�O�U���p�>lHu�8ӌ'A�c�)s��+�1�� 9,��r�z�OZQ@X.	�ZO�YUK�n���6Z^�W�jh�m�|%�O�|?`���mf�<+���(�>U ��\������5�#����#�	(jHk�:�������G�11���X�ϥ�IY�bj��_d٦VKO^���ԃ_�m���V���5�O�R��T�q��޿K���70�;��Ǔ��dQF �*�&q��ˌUo/1�/�	^�W��6��6���f{�z`e�솚�B�w�S�ԏ#U�؀��O��f"\1s�}�m��B��\)�s	f%9������*"�nn�P����ד��]h«�c;nEx���x�Z(/���e:��_�gHr Bh�A8-�i��f����H�i�?x�� t_AL��Qh�R�m�����;�9.�y�?6a�WVV/2�'''	�4��9�p����N�D2i�aN6]�e�A�e��@u���зn��S":��;��J��_t�$�9ƻ��Y�b�"V�o��Ytq�����J��G"����ӵ/$������}�w6�$�۲�`��,`��y����C�Mi�6 ����#�X���J�:����LN	�m��"�'>�٪������`��-+��)9��@r��--����"�!BJ�oװ���{�M���ƿ*e��'q3�o�Tɔ�_j��DH������QSV����	�HEhT`}]�q%0�p��,ezD#U��N:�3,.�0ګ� &���X?�d��=	2��F���:a�aEC^�M�,�Baw,�yoG��
C���+5�b���^^T��]`�>���1�l^"��:�#���烞L���O�aaaMVУ1��; ���Ы������U��+�*���m�J�b����ۛ���v���B��7��M'/��a�ނˏoj�$�EP����X�<��?3/~�i��x�*e'�hA���7>��;ɘ�/ �>*�v�Q@kͅ��"���T�����2"4N�D�!.g[���Y\D�	�\PJ�>z8K�:��1�m��1��19jU$"�FK�I]oJW�尿�B�}���QȆ(��@��w�vQ���n�V���pp:�0-Ӽ�P�\�I�˱�9|��5(�>Mz=n7[8ڮ�ɢU�>TB��Zh>�Ǒx���n"U����T����pg��ʧ!��es���Al��{kSX�����m��>5
.�oo�5:�\���*�;C)���FU�2���F��N4�4�_�*�ݮ�P�w ���Ꮣ��ü�4NF�����Ӻ<�/�,����-�<M���-Ւ����h�?��c!�Eؿ����A��]��7.r�f���sE��cge�l��LݫXӀ6ն�������^c�x><T�w��۾ͲD�ײ�J��ƖϬ4�`3(L�Z6�$��i��q+��("cNur4�r��s����	C/��u��W����g7���wa�m���}�e��d7��nV�)�H��;��$7���U��r�&��(B��*�VݎBs�"��Gq�Q��5>B�@�)R�i<��O�8�zPE�z�N��z��RJ���o����:��7���o�[GR�J�a�//!W��<�|Ɉ�[F=�v���`��y���Ո�K���T��>�A����σ)�_s5����T�~�#��Z1��C�c#����m0��8���s�ʔ6�"#Zg:�x'I�N��G�X%wiݯa�/`KK�F��Ր�Pn33�i���'7�\�O�%�}����m�ߺ#c�w��LoW�+uD���TO|�����1�!�C^����]�|q�$y�2�R�)�!b�)ck�ρ���l�@ӀdV����"�ݨOb�Q�T������!.���6�F�	�:��" Vq1���w#rG\�D�RFe<)C1���=<�+(�O��Yހ���b(3���tv}�W��nLG��Z�D��$n���G7��~�Ъ��Wad(�'N���U�N�q���[��$�w�q�K�O�4 7n9E6���RD�礲)�T����o]��I82on�i��������uw��ܾ���#{���(�������=k+D'�MXkDC��AAA*P���D�R����$��c��Y�o�$=�����Q<��𞊻V%��x���oN/���o�7�s�rЉ6��Ӆ�=�����|�7�AZ��q}�)]`� ��J��+��a�]E6��$
��ll~�9P=�w�&�B{�c�A%/� I��Y�9���M*�}����R@�.�
њ���>�^�Ϣ����M�'\�e�f�k��ߧ:ςF�Ń����$����6�{��xe9\��(W�9u�q�?1��������
�h�{��H8k�ө�����=E*�_m�g��	@��=[м��B$��e��^8'������`u�(���o�	4ayktM��ͥ�c���u�#d]���.]�u�������o��D4�0�	��Ƴ,ړ:�j��w�ȋ���[���My+9s�.6Í��>8鉟(`�z���N�.t�4���~��5�#u�\,���&�9 ˷7�������;�?O�$:7�6�K&��Q��ahc�j��@�d����YO[a+��EsO�ڞL���$t��,!�Q��?���
�q+T;�k�����7�r�,��
|��`��\0 ��5�<ܱGq,g�}ܕ�!Xi<5��o��������9������ڱ�hoˣ7S�_�㓍, &5jcE&Kaiྼ|���{�Xt9���}������9C�踩���Z*��	�N䬇���Q��>�"��B��޷���z�PjT"����ۉP4��~��Mx��}��#�[�B���#��l������ ��"�YǩD��wǣs�����=�ڄ�k���v��0@�(�zi�＝��qڜ���}ܬ|2�~�\��^�_ә��䌇�@ ��t�5�47t��ȞL
c"�����N/�K���3S���O#Kq��	�2�,����V�8/�/n1�7�&(H�T1���\�r�v���)Q�,�M�9�\�0k�ߊ2m���͘,�o�Q�Kd�� �l(�w_�1 ����о ��,���u��K9K�u����4��M�jv�����ͼ���t�E1K�-��2��-�G��\�˄��/-��Fŧ����$\�x�C{뮱��h!�]X�y�,��Ɉ�?�)�j_�D�c.O�LM6R�|��sՠA����@���ߛ�3�
4�y���H�ʄ�7[1~���o���"&n,ǡǳ�2��.��3�ۛ�O���Ԉ��A����!k:�VC�ۄ�2�gqJ�՞d�b�x�X tM�
� � .݀hy�='C�m{�z�2�ĸ�.bNc�� �P�ǳ���E�I���6��]��[Nq0J�$�՜L���i:-��	Z���7Yt�_�L�7��[��
Xq�k�WQZ��>S�2ReYBׯy$C%�3�'r�Aђ�^N����4T:��G ��H��I�qF5��&z�3���۫���4Q}7�I'��X�����yǒS-ܻ�SD���
����>�gC�ٞI2��~$���e |�[>g�O� ?'�b�j�A@�YY>a�k�
2������E �.�����N4j~L)	�S*�k���x�?��NY��|�g�=�b��٘
zb�4({���у���S�ǐ�#�-e鏳7LQv|�kX�FW""�j7j~�H�[�V�_��#�*�
�/ƴ'.Z:"��"��;�K1oUh����P��z����H��,Tm3�xX<�񔓫g}'i�:�#� �} vp��Ԩ.M���b��4�D�r��I��!�C�!���Ք��l�I�`$����JЅ�c�$�;���w�t=!�&](]����pk�O2��]�|�UR����>㔻ݛ�e��^Pq��V�#ş1~���ׯ?�2`��N�m���u��D�2��+�3-&%���PH�3�B!���:���$�����:�B�J=�s;jCk�b;�
��nu��3�J"Qe�F��%ŷm+��Y��%e5��Ȗ�dqj>k	r�B�vtl��g>I�i&v?��x�#�-�ŸH��j�R��[���A���u�Z���y�D��1rD�%4\�������Z���s%i�A�D���������"���BЩ÷�#8bADDTI�Dp�u

2��f�X����r�'	)�h@����&N��,����a�!GBah�3q_�|	<X�����T���m� ������^���[��z��
A�HGBI@�d�E�`�Gh�7X9<�\��@|U�=�$���8�[�cp�-�L�������cȏ$�)��?��c(�B�x1p�X>M"���d�`�w@��[2��,��S@�~..�0�1n0�� f#0A���v	�""�8`�s ��<�`�	@� )	oEZ��,�X��L���/!��Y�"v�G� 3a��9��� ��g(�A����$	?�&F�@$Wq��NC:�'.ů����(d��E�M�E�I���W&� ���ǎ�AQ�MC�95[�"m�}`@sڠ�9���ϗέ� �Ɨyv��|^��6s1��R� ?F�>�Z�<��lE}�o���������u�$��T�{> ���((BGk���=��q��)(&U�3�ܕ����W�j��p�Ȓ��P�BF����`T�� ��B*,=w�\w��W���t_�����T@|���Z��+(�s�̧����oK�"7R��A���������j>!�C�|�Ə;P�˻�Ԕ"�����t��p�R�� wU�?B4�8�-"u��� ����P~5���u�V�_R��Zi� q��]�'�z����Õ9{�!�������跶*�	�\lEo\�T���R��-����xV KU9Yy݈�cNp�w93������M1�s��V�Zk����j�[>8B"@��nNoh��9�9"��SJ�..��FڔW$Т ��䳜~R�ѢE��.�4��X4Jn��kw�3j��Q��_�����.���Ln����D]�9�Y�|X��kۿ�S�W o��nȀǃ��o�*�	��A#uӱ�m��{Cm�}'*U,D}���6����!��_!J��G�;�~�?���o�
���o>k�4��|r�����y�JӹkS�����C�\Xa	;`+ŷ�{,���?+v/�ꝟ��CFzn��%�
]�����&��]�H0W���~[�?��@��v��B���8���t��%ra�ƛl��N��јϩ+6ӊ�q����TP<���g"��Ôb�
���g��U"z��#�d��cv�$����E�����s#���~ˣ]���e��*Z�
�v�)��v�LQ6\1���z���(��	N�M.	��W7�vO�l���sFª��m�\��3��2��vD���R��	�1Cw�G���!��S���F�qf�u��Ҟc7��7�=>I�R�����;1Ϫ���s��F�#Ud��0ѥ��Sl_�zY�ͩ�����a��ӳ����"�/��S��݄�u��d�F�b���g������!����R30�,�JD�Ѫ&AqK7���� Z��z�Ă�V��fi)+#��:I�7d� �R�/��7 ����8�Wq�������nӞ�ܤtc��v��9GA�]�'��'N��������y�އ(E�غ�2�-�Ղ�����(`��G_�̌O}��=Kx4��d3rF��j�Q/��H��}���|^�̻[�`�T[a�f���r+!��F��a4�d��M)��|Dzmf"�*1�f�'��b�?�{�+v�x��j
p�h�D���G+��WǕ0�n=m?~=���J��b���ή!��h����z%����<|�l�_Y^$􎠼A�c��e����-��p֝����=���K�et�)�n�|u�k���Z�s!i����.�ѕ �p�W1�!xzb��C�=U�@AM��Y/��7 �-3b�o�M�D��8�n�%���ΊJ@�kf��� (�|�+-���(^�:�S7�zq7g�^��������'������ߎ����Y� Z�E*����j�����qz�|���Q��9f�ah(�����}C�5�u���d�=�_|]J�,�@pFZ�v�*�����F�(ٮ%e���S������K�ۮ���,����Dڈ{�{K>-
�,��
�;��ƍ�7}ܪ�+�d���!�"�X��X�����]��j�m諛>�*���kE���	̻���<h��~)�|M'z��>�<����x1�[f,{i��=�rГz��\�����Խu�����6��>C����t��f⪮;�-9�u{&�B���)ku�đ�4W*�=���I�h��j(�~zֵB;H�M���c���}���PQ1f��
�M,�-�Y&a1�(s�zO�z7%�ћ���Wu1{`Ӌ�×*V�v���ʍ�g�_ȔN<~�؝J���{)��ߙ�����Ek1%�'2��b�tE�~9�O,է��Y�~�vU=���h����[0¯��z�#{:��Q!۬>�&�_Ӟ_P�E!W<1L��ō��1~����̻��e�y�Ux�.�.��?P��x�"rϨ��me��Y��-��,#���й�2�z�5z)���z�6E�#��%mN�V�p�[�r{36���,��|��<�C�bPV���vs�������v?�I7�W9�k���%qX���O%�Mò�8&�fY���Oö�����6�߿B�x��B��0��gv�2$3��8�������8��7�.�)�(\g�BF��$G�e6o��۞��^�k-Z��5ý��%ݓ�"�'Q\�(Դ�q�v�M�*��(�\�Tx{U�e٨RFZ}�И"�hi��[?��B�����t��h�����B�q4�X��x�8"]j��6����<��?�a���>N�W 1rm҉j�.��0��#%s2�j�n�(��d1��b�9zD��l��:�n���c�1�������t������N齫{�yLݷˠ㊧�g�܎>k=��v�Ş17�(g�I��ê�v6wv����Gȶ���� �T�n8�+Vl�+���t��-�T���i�N>��?���]Z�*B8���m�ⅿ�ZϪ0����H�=�k���һ���l`�r��g��t����`��I��fA�VX����-�(o��r�c�dOl�#��dϛsU���
��^�����=��7�����z��֊vI�&�'��\
�Zm�i�K����)U�s�d��f�>&��3H�BL�)�A��ܐ��N�5h�▽�r��r��(�V,�v�]P�~k���w��� ���}!M �k����㛩�)ׂ耡Tc� [Ϝ���$uo?�&C��Ӄ��kv�¥�pX��ԉ*��j|]�QZPbJv�8�ZvQ��{��k9DG	K�L�t��˓�����E��.����	���P?%�2��4-�K4rQԪw�2��R�~�e��|�.��3|�2��뜫&�)X��M"D����rt-������e=-������?��>�	q�y�K�Ŵ�o��鸖3p&�/Ӥ/��\���I�i_�7D��d��ׄ�h�u�
��Jp�ĵ�N�N�� |���R�k��S�4\[-_&�U��pJ��������{$�O�~��AG,$)�Jܺ���4�F؉�U4E���L��Xby�V��������".aeʣ�P�ᚙO�=��=�0�?7���{2�?$�$�1uͼ%�=p�"i_���,/�V|Ye���d�FLw`�c�\ҶS����WR�K�XX�|�˪�S�r�r�`���;Ү���dX��Ln<[���XmnmՉ@_����a�:��!�}�ٽ��(<ff�*�g+�xo�,��K���ٱ�#�J��`�_l¨+����l��ڢ�
R���-�)A��LZʑ@��3u��N@��\LL^f&b���LP�~���Pt<����ߑ����������\���iG@3�QFz���_���(����EI(�U��j"��\�eˊ$�Rlw^V&c�VԖm]��6��/��<<^��M�n����U�1��%�����m���F^6nɘ�y�|��~�;BAE�f��3���[k�C�w������4��)6I@�1�筡FVy 7;��[N�"�7.�.-� �1���a99�CF�2/�KGJm�KU�j��m��9��h�ː�%{��Q�mO�\f/����]Yclȵ�5`�Nb��v:���ul?�����4u��pTK�KRaJ�:sF ����$̏�l�^���[{��6����5���[0�%ڿ��6gR�oo����{(���ܖ}�[���R7��y�Л��4Z���Ǭ�~@�����}�d���7�)W�n�`��C��6Ӕi�y��u2b��H��(�1�	1.o��Q#	=P�,�E$�B/-QJԥ�*s��d��:?-sEr	/u���ڢ��w(z�qAYB%f���v�;���q���0�����7Y���3I��e킢D�����U7�`G�]��)2��j�{�W��/��P�`ꔲ�n�a�M:I��JH��-n�:4�������}�H���ܭ(��i�x�H����^+�݅>%�3�E;�k�&�|P�l��~�܎� )��M�������JWŉq�"�e[���{�v�����a`�� [Q�tģ(]�G��FB\��$��@v�ue_�
��$o���EQ�ǜiv	�eZA5'�Fw��~R������\���e-l,��
���}-���:��d�JXD'�<4�
�?_h{fO�U�Aź%��6PU��'�O0$դ��_+�'|�HJ�ms!�W4��C{X�<��wb��rͫz��O�|�A�fv�A� ����=;�ߋ��rͲ������rhfD������x�Ҍ�[7�vQ�7�`?�'(2o?KW�8�Re͓G�D˘�f"$D�&��tbE(¾R?�^C��m��v:�q��Ī����ϯ�ܗ���p��)�t�J��{�R�d�Pb��$�-�T9��kyP^7xKW Hu������ ���>�.m�>�hf(fI-�)RT�)&uj�{}1�w���4C�B�#8l�u8��;�E�Tg�+D�\(N�Y(c�^��98sd�d�����ȡ�@E�+@GdڗBsa���X�5dH�&��>���������i��$"RC�7Эڎ_�,�h&����+^4�1S�F�Aa�h
�7P^�2������0l����7c���D@(�]+��qC�P����������$Jo�$Ni��5*�ɣ�tb�8�T���~��4��j�EoĬ-q��r:��6ndE�E*(�J���\���������q�:�8ј���բ��b�8tAZ>�����~ևH�������ZKn�O=�l���Ox�Y��Q�4F��Z���e��Eڄ���^FA�ݽK�1m��u��m�x������������w؃F���;T(U�b���`jb��9b�*�ub���[k��*zDJ����L&�3����7�W����U#'�Ǔ�l�m8�9����)�*���3����*�k��}"�	tֺ+I)��p<�i����]گ��)׼?�#J��/�Ď� �i���g�k� �Ӌ�v��`�cC!Ɩ\�eO��Us#��ΝQL,�\��Q��1U��n�nYz�x�&SV���ߵ�{@S �~~JN{k|���9��?S�Bp���]�M"�5���zRv�:U<'��r���j�F|��܍f��P��}�Sgn*R�~��N ��[�V����mH�R�`ݽ�@��x0f&|B�W��Mo��H�J��B	�����%�*�����}�;��R�+��#��)�j��H���2l��+K�S�ٔ�������.�f���ȹƘ�	��W�%�H>l�\���kq�Z�gȨ����e�X��z�t�����_v��|�{*jC�� �,�ߍjfC5��a��:j���y!�*�bbU1���Sk!Q�-������ƴ�hɩN�fS����@XNċ�`�ô�XDt!�J��(%�4G���ZGo}�,v��I<�Q�uaz@鐔��2��;f��ӛ���N�:�8Iz�Z�"�mGW'�(�r5Hr�lV
4 �բ�%N4bA���#���?��IB&�6H��X���n��wy���î� ����$!G_��}Y`�(���"z<̒����P���[W�m�ۋ�1}"8��q���@9�S�%�	�&B��SN�l��i�-�Y"��D6̱������ɻ���_�n�?`4���P����Sέ���C��K�a���](�v�R�		�E��V�_�*CG��юֱ��|�Y=�(a�����E�6�y�8$����l�5���2�HtLKvQpZz0{��d#n���h\�Q�̓[Q���2{0�����ɲl�@=��` ��dԶzS@%�P�A���D�!i=H5>����A<8���*C�mx2��Dє�D����+Њ��(��;�x6J�܋�.)|!Z��?�G��p/@Z��bL� A�K��	�	:�|\(`$���u��fL_d��X	1'&TJ"�)P9Ef�\d��t����y���ʻs������k�s��b��đ+n��rB�58��GS���b��L�^�.TIzĭ�fi+��$$~�nB������2O������n��en8N��).�cf�J)�W��{Y�}��x�d�5�(�"SZh������5G}8�~7�\~�	^�`W�)�����O+���C�Ӯ���{
q�ڠ�ωF�:"�N>��a�R�+�R��ն�����L/^+�!�Z�~�
�I����D����¦�f���~�k�K�{=;�`cz����e���
��U!&�*�`��}<�c����W�0D<y�3�X*@���z'hyBBf�� 3����ࠇ���:|�օ�.��K��e1��
����}Cn�#6�^Cr.PE��)!�D̯q����G}��Zg�����<�w*�����t����Y_�R9ݺ	ǜ�}FN�3��ǚ#�?�א�><��N����9�cy ���I�'�01��(����g�w[;���S����aJ���g��=�O絮�L[3;֜��^QB̬�1-�̭3A��XF�dE�;�Ui]�g����:u������Ev�+�zI��Z�JM�R��FZي&]�<̞���FI�&����ǟؑ�ڠ��1v,&�@��4��ȾT�x�)SF�:Y[%⠇ml��\���]��H�3�2�G�%��\Y�:0��L��N8���m���3K�j�}��Yc`���̞�+j��֙/��E��H�Ӽ��0g�=U�c;cM����NE�MF�����G6@�-NFF����/�����g�*ӡ#^�RN��Kl��DEE!���Zߖ�|���	�ֲծ��,	gJ2���ɏ)�L�U\ω�jq>�]��!;�3Qo𸲭���VѺy;c{��=4镻��T���>��߾���x$��Lr�,St (��|�O0�Ɲ.�S*�'�gi�~|@���*�}m��V�|^]V�Em��������v������cGE[�<V;X�Ukj�6"Ù��߿�JLR;�y��^�1��C��kGOh��L�Z$Z�M)�ϓ	��)�&Eү_ݷeS�ݭɋ_�,�s*H���Z����C���2��mN�hP@g��AX�a��X�����je�3侒!ݙ�R.\ޠe�@��ɺ�Ao�f�D��p�L�`e�>uN$�a���p�'��#O_*��V;�~�Lc��GP���m�;��$���8d>�FT�����$�0?H�����|%Ĳ����B������%�k�?�E]�2;R�W=�C�9ԡ�`
1[6�'n����﵍@��v��8r'��%M�g�'~�u���W,���-FQʢ���ıy&|޿lR@����~����Je��w/�}������4�I 	=�R�l�/��|Q��w�[^b�����||�V���UM�@ڶFT����7Uc�i��W�O!�(�޼�S���'�����7�s��f,���b��U��GuE��޸��	������_T�8�	ь_�y��_S���Lq�"�G��h�4Κ�®��!��*�؁�z1f?�(Х����������+ �:G�������㙶8U{y�ਔ͈C~��%��O���h�����ւ�/� s���5Afe�B�J���M��l��@�������'-(�PZ6�� �yOOc����/%iC�ү9춧�.ؐG��̨��`�M>��_^�6��%�3�q]�;�3\���6��d���~�#V���Ћymh��6K#q�����C��Í!$�?u���"5~��Rm�G�k�m��'t��zJ)HN�HW{<�u�Ax=G'�ʇ|�}tt�\�􋒲���NU�bПN�K ~��g��)L���I�˫0�i�ˁxG�R�܊gϾI��}D�F��aK`����=�0g�U���f�2�)&~��c�IԻD�'��|ֈ��Uoo~7���c ����(�/d��H���6+1��^U�@F4���/d*X5�d<M����Xm��dbn�)��TY�s�r���8ؘ���i��L��X��x|(�uj��g���v�q�WYܗ��-1ډY�D�}�1)j`�L�}q|�VO+���wX�k���#�s�N��&�Z�o�^�ĥ_I�� ��w���y@Ũ.�]Cs�:���a���T�g6��ps�|2��c���	��7��L�5VH�E�1E���~���D3��4���`/K�7��#�T��H*u��n8Wm�~��SQi�_6�_{z�j�7X���RiĿ�9.=rM,̭��\�Ǒ]�f\�(t'R��ė���P���V"�����Zz��T��N�2� ������7�e���wbV�@�_��0|��e}a��oVs���ܓILoYa��7�f��&y�W��L�|,�E1t :�k��i�CD��Y4t����"�\�$����<T������9��:�d�uM�L��ZF��R�Q�l!݀����P�?���N�}�0��L;��=0tL\!��^I��'��(���<%2��V�t,�h�B��Mt@���$�|gý_P�*�>S�{�"�x�߬��QT�V=sTK-ê"{�16IG*%��;ʞ�R�����ݹw��<_w��=����c|B)j�0�X���A�3���"k�s��Ѥf$[�c\zrso�[�F�rXy
����"�����x��.�������h����O.!n�����'喭��-E��K��8�<��̱N{0�ge��<S1ϭI,iB����BOt?���.Dwt��+���|�{'��_iؔ�w�����Mga*
V�\59����"n���3k����)�#}H�{h�h^ۄEr��< �n(b��{L�{zDz��j)d׋����mVqo�/-$n����}��D[I>*���2e>@p;���@�7�؆�'�H����g*��t
S���i��f�Aڽ���� �?g����_䝽�E<�hO�IۑؓM�V��d��lK���b0�a�_�bF�W�`�Ա2}����ej1@[���X`�B�¹
g��==q(�)"���I�{�r5貞�4vp���s��h�W_>V��ڷ�����hؚ�����MBD���{�1��y��O��U|�]���	c#٧�8��Cp�dC�E����Rve3���ձ�r�5�4n蘭���?���#-2�w�z�祣��i���P���բx���p�Z�}�t)��(>���'Anǆ� ��"��o0n�L�g�dr�R��b�$fн�$_���N��(	�S���5glc�^/az]*+�z���҂�k���	/[��cPC#�2)�Ԛjv�YXy�mC���ʛ�����������PG`v��AM�$��qar��d����h���ؖ��5QiLZ=�Tn��L��K�#(�ǣ���:g�� &�B�rx|���V�=�}��*��i�7v�����`o�t�ì�%&�j�
mu�x�<�M,�)�QhR(��p����[g*.�j���M�m5|1�A��Q?�����y�ޱ���c#�;TJ}U1�O����]��#��eI"5�%�}��:��:�Ӝ2u�����q�R�">)x�҉�9�����s��a���7`eI5:�88�+Tz�v.b1.�Rk��)}�ݧ^Z1`�����.��Y�n��3�8I��e�� �]`�N⍂\�	=����m��#��%k����y�;o���q�?L%g�EYik3�׆\dk(E�H�:w&��$o���C���u.N����:�E/�M,89��u:���K���m'�����h�9&M����2*j�د�����Y����	�&kd%pC6����]_q�"|�'��A��1we{�
�_�+"�������1�^��6��؊�,�W|.j����;�g�t]��;�m��c۶ӱm۶m���8w����>���h�k��uUͪ�Uc�0f�j�Գ�++��¦������|�B�0��1����Qx5����{�RV%�-�컜.�m��I�PL���ga���?v�b�8�jE괈����v�2ҙ�̻�����l���N��������Z��4s�#�~+eU�f����H(UK�5�U���u>��Yr̈Q�����R�$�`�ik������6��v����T���|���bQ'����i:0	���f�7��Y���Kic�-iW���Z(������g�J�6���e#7���c�Ob]- ʔ�N���2�兛�f�j;3�*�`�d��d�]���b/P��BH�:�qo�O��2���w��[1ܺ9ӊ�9v؝{���^r��4��x�oBš>��A�%YX�ϕ��uTu���M��O�f�6��,��'��/*J���'� ?ENt�
.`�[1�N�_\En#~�$���t���s�q�E�g-�Օx�� �7ѫTt��|I�R�u��DG-�s�<Tr��vue�x��69�#J�6�+��n����	0}���@�德!�>�E~/����A�M��.�\�*>(pm��8����Y���GC����U���+��rii_MЎGx�꤈��Pȝ���6��%D�����O�'��MY�G��������lT���6�/�����J:έ��*8o%@`y�6����5��U�QʢQ��;���v�]�6��� �m'y�,�Fmt�D�{�y��)R��CDYH�m��DAD���HG��C�Zrel�&^Eq�������nY�z�|����Z����a��WK
�d%ɏ��2/��H���Hȼ��
���(ִ�DGt\T�H���ge�@���,��o��0WM|�q>�y�D45��H��)���I���zrR��&Rj�ABيI���ӂ�H�+�Αą�_7|�x���e�e��o#UZ���EY���֢�U�w��i��J�z�,Lc�B'a��ݩ�j���꽗&xj:�3&Ԣ��=����E��"��Ɇ�����.�u�j��[�1����>�c��?K�ψ�_�rt!U�7ߵ�V�����?d�$e6D�����[C�.�6%�A��I[�v�zA�N�r�Sy�����5|�������J��Q}��&���(g��<����
��j{d�U��J���Fk�Z��ݗ��{uh.��e����N���վ:��|F�h4�R@�X1c�i	|����A�j*�@f�����w!KzUx�
��燽6WsD�ۓ��j�@�^G�A��sX�4�ox���1�{?=���݆LG^��Й�4H??�^I�T/����2��Ad�1�%�/�p�e��[�����"�]�Ґ�ز�h�<涷/���y���$#�h�x�3�_F�hѦ��}4�wha]�a9�bxI;����q�D�,�c��}��=/P}. �Ӎ�q��p��Y�l�������=��T�S��������gS�/�n��
�P���~�����N(<"k�����Zɔ�	06VC���V����K%�򻴲|�z��C�^���*�K�e�g5�����o���y�L�����'8���a�搑 ~h�	_�CN�(�ص��� ɸ��)�U$���?�	#����e�I���p��P�E�
-���Y�t�W*u[]o���-ng�u`����%�����=����cF$l0�&v&�3u;=��GȋeG��5�򈗺��n�ԕ����"�L�T�Mq`�^��iZ�j���"�+���p�T�k)	���Rz	��g�o'���_~"���;�@Ȑ��k�F�ЧŜ
�,ҍ�L/x��h!�@�D��⤫�!�@!d��B\���AQ1q43)86�mi�.��
�:v�7���r��*Vg�T��_M�@��gV��z����ە�o�b�S�l������ k�g�KAڒO�;�jyY��)�x���{��A�p�T�ϯ��J�Q����[��J!d;~>L|[c*eG�<��#4� �(#��U!���x��W��j��j,R��罃ꥅ�'���`�+�Đ+,�{W6���G#7���_'����L!�GH���$
nA����"�}+u���~|����q������|'�IXz�y,FrC�e>E��P�G!���'�k>Ɛ�gʸ�NR6A����ϰ��`�W���4%�����3g����#����06/���@���.y2�؄�$�M�x�L2�?��2�&�$�Z�\�S���&�5i�&�Zc�U��`{Y%�!PN��PSl{Y�6K���!1��/S3|�����P����
�����I���G��0nTW�_��Z-t6ꐈ�=.�{[U��V��P���4w�1��5EÑy��Q*0�Cicҫ�v�����a�X���N� ~Ia�G�K�tx���٢,�Va�%���i���0���Ős�!��N���J�ZQ��Q�e\*o�9�)u��p�'��J��T� ��ɤI��jѱ��(���a�a�������!�~�tLA6*���ݚM�h\�,g��ߔƙ���2�ϑhV��g*��:V��"�K`����V�X~+���:;���M����:]��<�-U�q<O����hw����/
���%��o��(%�WKv���4Wtjy��ر�|죻8�E;v��
��)L��.����_�_��~![c!�̄�#[���7�K�.�RE&	�CHƔ`[H�.�L�O��L��Ib��(I��!��/~^c�asl�6G��f�v�z>�|ݪ3)����}�"A7��S�����mU�Z�Ҙ.�@c�1���%�|��q��f�MU#��a"��ӣ\�6t����X��3��~�cS��E@�X���+�PG7W�x�`��͕n��#�ۣ��7p��PP�tb�ʍ�s�}���tb��"���a]h̕�%���;�&�nl�}]���dc�^�wPI^`���X(k����^�e� ��*�l�����E �8�K���{�Z��ȅ���@u\�T�g�.Q9k�L���Ӫ�+ěԀ�y�����~Lb�$e]��@��+t̃\��Ĉ����u�Ɓ��J�@��"j���p��d���F���l9yA8��a��D�G�Gk��ʒ��z�>�ؔ��9�C��~���{���n�d����(��6�t����o�uQe��:���Ľ��h��	��1�%o��J=
F�|���cǯ$ζ����S�ϼm��梕1�I-?�n
����?���u��Y~��rm��������h
W�%^k�v�'f�M�ɀ��;��6�z��ᒭ�AC����J��������(z��}�O��F��f��.�e�=2R�Z2��yT�d���"��)��x[��ǯxGр����ج�\���`6�� j�f�΀KF;;)�/FlV{��M�zHt%�ź�e>�:Ē�1||�ٌ��E {�.[w�����[%��RR�2�^S�P��Qzj�rߑ��Ġ|9$�:|��r�A	7�8\���	�r��.��d��^���}����w�줖O¿������b��/� ��p��z��\qYD�o-Q��78��,��Ǫϐ�)�D]� �gWݾl�@tܤ����z]�#[����� ���s���t�:2�2X0�Ov����� �k�mn^�y��g1��@�Á10�8�`��oMw˯/�;�hʡ��d��g�B�&]àQ�V:�YO��u��^��֏{{�OoA���y�A�]ة-p(Ao�瓞��j�V����m�(�]��0�<NJz~#������J��;^������G�`W2�8��OCV�L� �q"���Rn���@���$��;y:)��c<c��f��b��@�)-�v��.ޡ�{R#��iC%�����BY���T�����3<�~��(bX?����8E�^�lw�����-��@$?K���������v��u/���F�� �g�.�<R�av�j�������'KG5`P]ؖ'ʭC� �]�ͥ�G�[�v�{G�/M�6�`EC����As���Qܓ�������e�'��_%���`�KZj`O�Z3Ĕ�l&ŧK�U`+h2�-��}����u��e��e)f��k��(Wc!��O�10�q��u�<����eνm��I	iz�ɺ��{��s����J��P���#�wldS�^���#Z~����f��N���$��F��ZǕ���Ĩ�2�Lі��.<Ώ��|X$���EϢ��_3V�VI���Rp�*��A�v�����3���|�L��Z�ϥ�A9W�ҟ�l�������~���?H
59��;����7��	1��ll*4"��:0y�0�M��K�b{&t�H��V^��3@���wr%�v)93��E��p@���BO�K��?�:<2������7�P>�|o{~;پ_uB�U�;ݚ�����3�0)w`���:U�1�(�n&U]�̞�{�֡��
_�O�_al���XN����bA��k�8��L,I��/'��c�gK�ƽ���q��G�ķ��ȱ�BP�ڋ�������S��^�;"s��*�f�jf~��v>��j����p��QQ"+v��c0�3;�2���ñ�hI��&4L���&JaM�X�
A`.:_*�6��$'+�k�?�n+�5�:F%j~�'�R���b �A��!�3�F�Lk>L<)׆�u�T=�UEɎA��lF^N992�u�ߦh'Ɇ=��P����&rUN�{^�b���Ĩ��B���������"�6��x�l����� �|��������z.�����Z~��B"'�P��<��,�H��O�1Gg3.N�j�����xA��L��Js��y� RIP7�X4߅�0{ҙ�ԗ�YE�&4�˯��e}��x��i�C�P�o2ؤ�&�&�"\�����+�A��^�>�').���L�����9���+�C.971�N+�yP���Pr�j�ڒ��K/DxCG¯_��a�Bm�9*�ܧ�|�$���'����u���Bx��x�x��&T;^�����z\��
J`m�H���x[��$��//~چ��B��A�<qM�����a��zV�Ǫ��y�,�PAE�*f��í���mK�{��\��	D�hVvW��l�M,�ʱ$Eؿ*ks|t�$k�����L*�Cyi�5⮈#&
L�Nj��$ɰ8N�$K��4��q%�c����`ol�Z�t�dU��&�^�UT�>~KU��x����WΛ6�]��l�#�h�g�q�&>�1Z����X1��F���D�1�e���K/�^Z�3r?ÉD��t���8�+��%TK��_�%�i]��1D����B�G����~^Õnk���/�u8d����ƙ^�,�]��O��4܆�ZP.��� �}Y��c�9՘aLbka���=���=��H���Sq��\)�,Us\j����j�hҢ�ST������Z~����v�O�9J��������0آ����N�I��3���?V�tMJ.Wn�rE���p��)-O���}ا�9��R*B5�%hdiPt��*�(d�]��d���\g*����^ޯWL��z �ﺱXcE/c��M1cs�y��7�z�9�x�[�߅$�J��?�e����[�:�n��g�
ozzs��{���+��]%E��yN���)�	�8~�^-���A)Ɖ���V��P���z�9�IF�S1�O����&�]���c����gTd:�#>w��e�?,#��(��"LM�3R���O�����x�O�v`E"Q�u��BPp]��RN�_�&CJ���� ����Pf��C��`�{<NIe[�=S�5E0;�C��!K=ET���[^��'�z��J�dNyv}�Ev*��Q�F�b�}9�x����y���^)��$��j�8K�!'u}9�lB��o����@��S1��z��x4��:*˜�bp�`�c��H!릵V#"�����8�/2�s�%�ʦ��jp%`�#/���"���͢�������҂N�X J��W��;xJ#���0�T�\>{|�L�?r~�nr�LE�)��JN����A%(�˩���IKu���`����fN�lq���P�BO,sC������h�6�)��%uO���O��g9 ��
���9R�!���Y������E\�w��I8�4d�l-�wp���
�Pk֝��_�"��&D3����w��d7��Ta8s�χ	����>���9J�#�É(x�E��aD[�̖�H�[cH����B�����y��T�iI.�ă��ײU��O�f�(�v\��aR	xeVV*���.Mנ8�?����b�'H��%{�fo5V�
qE�N=,
UP�����rY]1CC>��CO(�VS�S��������V�D�W�'�M}�W�{�t�Q�@��O>��Ԧ����� mMU�uڭcX�
3��
OW�8��9�&O�%,0\E��?��@��8��~v9f�~B'u�SOf�����έ����I��8b������IB$[:)�Ɛ���^U?��}#�����efxi�;	'[�eӰ|�y�&�@��&g�]�m��Y� O�!y\��N���^&��˵�t��cEȎ)S��˾��CUJ^���`����ۛ$v��ApJ"G&�W���O�p)�O��Z��4��2����TU�o�����w
��1�Yq�(M��H��o��I,�7>�w7��A�������Xb��d��kH��s�}����$�Dۋ�����_�(ƿ��h�}���R�?\�_f��bzM&��,4��y����T���8�ا���H�����,G�XO�f7c�`�����on��%\��w4(Iٜ��&!�}��W��1�9���>*��z���'�(���3|a�:y��E,���R�G�d֣�,4�j��߽�W�yS��B�#�m��^��^vwۚqb��(�M=7�Zip90s��4���!��#�C���a�L��lo�sK3@/�θ�=30�ɭ~�+�����ӄF,)-�J��]�6�<�5�����$57���!��c��?���FaK,�P\ԛ���ꓩ�6!���m���;�NtnZ
;nѸɆŷO�m[fn-�$�x�c�8�)ت��˭_�o��B�4��a���]��QO$���@�:�i��!?�wP(��'M˔|?����@�K8PЅ+{TH��
��~�VU��j�9sY����O {dJ禾J�@�$��K%J����v.�����گ���v���������c4��d�� f��i:߀dz�i�u��}�+��2����Sy���-f�t(�����\鍰XpvC���|�W���[��z��,��_?;�;����h��h?�9J�L��71��i�e��i�?���[	O<>�.����)&�G?=������Z*�B�\ɰ��㌅�Z�ie��V��(cn���s>P`I����=��CHX�>���_Ic|��ܥ�H����;��7�J�(t;e^�\Ni�j�.9"?fHe��=�|oa�7�$ؿ�t������X�����������.�a��0�+��Ҷ��E��;�?0�N�����N�xHKBh����_%I���2��C62��1������͋qETI����"��Bt����!#A&h��]�+�x��*���#��~�;�,�8�	S�X�^l��N��!�?�M�@�V8�MySS0��VoesV6��Z
7��|�8?�Wt��#���H��շ�f�db.P��T�nsȏ�3A/<g���ʇ Z0u�s���Rdu�{��i	DS	�Q���S�>�z��|z���Qo�S��4Y��-��D��erǮ�>�{Le�>�}�Q�R�P�>R��&	���v�I<�o.���1L����~Wy��s.Z`�Z�
z�����
��5d���n-�}�-|E�j!(�nD!DC���H�!�)�*�jPS�)�O���"�|ຟ����[9�tv���:�.Yk_���D&R��m�ȉB�B���Cr`�]��t�ᾰ�_�	�Í��gWk:T�(���8�
��F[I]�f7���d�o�R�$Ŗ��Eau�c0m}�Y��7ٴRP�W��Y����o#�w�+M8��$��<��@:{N�`�å�KXI�81Qw��6��-�P4�WcfF�j|�]����&;��s��j��N�u��7!Mn���@f���{��Q���(����7�W�7w�N��`Ö�jڣ����:�v��n�G�:������U��`/���.D�Y���H�ۣ�^=�_�`b����PҰ��j��5��{�e>�e	@ l�}�A�q��g��]�褧�@ݥ:ڋ�O��(7(�P�%���D��x��d{�M,t���T�FP3ڛ
�4SzE�2��Iw�#���X[�D.ӳt��GG&4T�ϔG/f|H������������M�����	-G��c;�͝�^s�>M��KQ�9C�#0�gF4*����^�E(/�E8�Y)�JJyVf�4[����'���sI@�U��p�=eL��t��Tz�z����U�!K�Ňi8�T��׵hc�Y�Ӕ��[����UQ̲�0o�����HE��i}�s_B�� h��G���-�'�����"a���"�uy���J:�8�~���oql��m�~т����^��)q1���+^�����YjWV�7r�JK����ؿǕJ�J���L�j���a��;,Xگ+� `"�}u��7�}��!Vs�秉h�O���O橩����&��Ҡv�Gw�׵�Gr,Je���3� ��K���N�F�_��P�����[��n��u�8"��1��
� ��0�P��S��ZAb�+p"�@��ϖ�>�R=�I�E�&��ԭ���dw]~[��[v@���ވ&3�AS*�Q �`��l���.40b?a(����x�G0a�ްd];��<L�	>�-.W�Ls@��_�����B���B\���9�8#�M�8��R@�]�<�cM�$�H�N���lkL_�x\m��>4�9?��ωk(%-�ND]+���uz���'�<�i�����Y�D����Ւ?-T�4��fNO>��*K�N�9W���UE_ޣl�0�N~�U]�P g���e|6=Td༷�=����^�����RA�@��Gt���*�����ݾ�/�f�E�a̫ k0I�����xh2X�r]��o��Y����0�4Q��Vt����AP�_7Q�Î�or(�*�zr0L�|�"58y|��\�k� 83q�g�D2M�w�!�ڪeR�]
�!\;i����U��.ے�O�LC�n�J�A@��D�U%̯٥���Q�a���E���K�$*�}��nPlk���2l�g2�Ûd
����ϔC.�b��T������h�wT@j�7���5>V�ĩM�D.�f�|�u�.�C�3P��$�q"~���[?����ר�2�4>�:vP��IcX�`1�ӏ�����ײ#�
�u@��1H�p�T�������ٓY��ߞ��}��n"��X[9��PU/zo[����G ��XE*�R�7�������QvsY��k󧜈&�\��g�p���j,y��Rq��jЅ���\ǎ��l�?<rGc����-@��éj�(�<�I�k�h��c��|az��q���m����Ғ|�ŧ���Hl-�5I��>z�	���*�^ef����6½���;��R�2�_�����ͷt؄m,���/�UMi���4�͖	;��6�'A>w�y�?^-p�EA�p��o�nE!��>�8c��u�}�����M��*�||���o�1��#�5&P�4���ڑ�,&,�G�0ƾ��mK�!���Z�����w�AIɉRy�9c׵]:�Ƴv9�%�в�>5�Q@��5(��'�[45	��R�KHՋr wޅ��w�:GL�B<�b
~s��=���˂�jB6�a�i}E�:�cH��]	k����?��VL�&��[6�"��H^J�C%�@,�q����kb�9�M#�����6	�^�D�z�+�Z!�4�I�~�Mu�k�Zx��..��GE���W沧wx'+��\9��-Q)�\�������)�ȂE�҂�Ѵ�fu\<>��^0��ww�!%Kŉ~�UI_��e��aRSN��b�k�*'gbk[��$I+�~Nh�ڋ�B<�6a
���`	'��I�.���A����b��Xj8:���٬��sj�kuS�o���]�c^�V
g9[�s���b�Fނ�	�Z��O`��]�ΠE�)�P�U~������	4��8/EI?���|\\\<�DEE��pчh@��V�*붏����Hj��ш+
�k�_�,bHn�7���w���܅Hh(:�y����2D��]���#ό@QK��a�)�|b+���K|Q9��7��o�r�o$£��ap~�(�_��߇)�kh�`P����n����D�J������r:#���-��b�KgHR��˷�XK�<�%��M9������7A"��o��te�g<����	�GֲR�X�޳k�2G���l�K�j������)~�I+Ot4w�ÉT4����r�D�BV��o��IN�6���_�l�ʆ�y99ق*�#�v���r >�L���SrT��\uQ%6�Fޤ,��� ,d�[�`a�+��s��A�Gq��5�R�f��X�&�{<����y�$�X��{�D��.��r�#�f���V�S?��ɶ1'<ߏ�9�� @�����XX��\�/ %�C�8x2�qݜ�#�TSW0!��QgD�)�}��w�(�װ�qB��g����r�t�%C����Ln���{H��ыR�b/#b��stŎ]�^�54�P��/X�TR�Cj��$�����Ȱ&�'q�S9*��"�R�d��|��N���$/(�>�	h�4Cܘ`WQ�Y�=�63��{3ĸ�� ����=	�����V�urFc��M���2! �5�G�Qά�v(��Fc�;I���wsty��E�������J��B �5StQM�N#���\�v�O���"+������^&��v�ʊ]�_{ns6�[t:�;��U��52Ƽ�I�;$�ƅ���Ky����?9-S�k"A`��X���O����:Y��I�ȳ�G(���/2�t}tەΒ�q�� F� <Mb�W�it������f�:������Z�g@������������oh.z���@�?��|�x[�8*T�Y��ެj�ykƨX�L%�F'��Ea��&[O{|nq��S����t��1�����Qg/�-e܈B�[� ��'W6-*�M�(Q�'���[2���X/s�a�
�d��H;�KX�v��K`�[�U��a"ݖ�꧱4gh(�;k�4�a��=C�@-Hb}6�=����f=2IT��� tPK�ż�9z1H��R@��Rt~��ٍ�����I���>`g���t��k�@#2_ZFzW�k/�S���`���0�/2�����]���ͦO�t�cp�:�vGa
�2'KL���]��@=!��4��� �D[��J����d�W���k2�c��Z�.�.�w���x?c�FP���c��=uݚ�@ ���	/���z�=����RL�c�`�\ZlB`�$�����#���4v�av� ��4���F� �U�2����~*��߬�qw
��S��������G�G˺�[C�
I������Ե��e#G�j�B��4�Biy? J���쪓j������3��i1��pK��(ҋ�o�lA���TG+wʢ�-[�D��ް���,���]s4�>Z�D� ��j#릊���P�c�v����d�JU�a�:���� �6[��"��bs�UPu���׾q��|����1�41޷��#Vƨ��L��M�N�.��L�A{�ƴ'�������2m�z����Sn���m^UV��.	ZrI�#����)���p�tn��O?{X���_�{�x�&�Y�pߧ�xn��h*�2EJ��!W�.�ϧ��;`���������6ӵ�4�o����C�Q�Qi����[w�GN�"�J�oPX�n��<R�ЮM=o!��wɀZ����>M�(VN���J����4�5�K��;�4�cP���\ A aЄ�ŃϞ�d]&�/�{ϩ�����n�&S�t�fHs@���ء����B�a�3��ӜT3�Vx�:	Fk:"3�������=]���bM��xw��;����ț%����"�b�>�p=D����{��Q����{T�ѐ��?�f�	w�??ZgHqv8s��9_}F8�6�Q�jO�;~�F�:j���j��s� ��joΟLc%����כ|"u����2l�[5R�!C4(ĥ{o| A�1����?�f�5FhS��IEC�Q��k��DBy|��2�LBC�6�£fv|�pЬ��ʰ́�7u�@����f����� �^�Ƚ��LK�D��5�B"=�h�����}o�n���Q�
 �i�����&R�#ѫ��S o&��q��.N��w���F� ��&׭�=d��I�drd)���(�g�r��:z�Y������I4��!# �䲃���P���_�x��[���e
k����A�X\§�h"�������U�Ǐa)���Hg�D��K7^�]2K���)(Jm��AF�
��G?���ұ�6����K>��e�j�R�����}Nqg۵P!����x�j�dXCb�E��N�}��%>���*���RU(\�O5�����h�O]`�
���2�
�06��{����f�]7�Z�I�$����g7/��I%����>ٽn?_�I��+�mo�����vb�ߎc6�߿��P�w������Ei[z�L����w���%�F�wYU�x��@�=X�L;�E�V�Ɯ� � ĕ��2wP���V�(^^@�.s�<�n�Zy'�sխ]
���c,@o2�����]��
ԯ��=�!�4�šX��R��Y�sօ�MJ���#OGFiԉ�"��dҖA<5k����nn�d�A��;��ܢ����7�����vA.�#�Z�)��DmĎ��j���51y{��j�B�)���_đpG��:I
�KhW#0Ó]��D"������)A�0h2T�@�TA��)��5X)�Kh�ھ��Y���PeZ~�IּKu�7�pQ<�N0r�L��а��@մ���5.�Wr��>	�|쒐�1~�R�NO��S�I�����8�P&_�7�T�r�H�"�P�OUr����M���j9�	ݮ�f�a�w��dBM�k��^BVXR��]��|$=��=��C2�ޔq�fF�G��Ѕ�(Na���Ll��"�H֚��!����
Qg?Z_�-I��dn����`��+���	�{A^f�D+�(o���ټ�!Y�O�%E,��@;�<���$�׊6Á�|M�wvކ��HJ���]���K���c�$��p��oc
}?�BChш���#����������1�����q�
Z�4[�
M�A/Ys(哋��\��]^p$����L�_��yC2q��P�8$��f����C 'g5��@�|����w}��A!Di�x��8�&j,��5�D�λ ᳧�7R�J>D����&���7qQQ��F͑7Wh�Um�Q���5K�̮�i-V��]�K���K`�8S1)^~����]yD�γfn��hA}PCT�l�����1����L��۩�o������ֵ�3�ի���s���_	�{���]�?G�sB���O���➽e��ѤÁB��wJ����8�G�3_�_F7����p��&�`&��5F�K���ɧ���,����9b����4���T���m�V��-`��7��:Z��P���-�ž��A��O�K�3��e��}Aso^��bh"aM��ғK{"o�J��H''!r�8����7`�I4C٣�m��?@��no���Dy�q�.1�>���d�:k��U.���6�����9  +
f:�~Jwo��1	��A$ΰK�Ե���D:Ju]l��4�P&�����L�5�L.T`laZ6�֌�)��r�"e�}�*��]��J��eP���G�d����H8#�0l"��b�v�&��6�6��Q~�E��"be_Q�=$6��ܫߍ�X�����⪬��b��������]H����Uc���f0(;��r�=�[���=i|�1��`۠������)5	����MAn�$
�X^V�v{sƼ�Z����$�Vߺ�Ic,�49d�hnNFECS�x �ə+$�(}���>���r��e���v����+�WX�L��VTSh�{G�o�!p�N`��V*-�ƺ�D�Ba�tP�{{�d{��+*�����Lo$t� q��t�3[�uZ$��e�)ʼ�}3����%$�5%½�p�P����~�q�檵�i5?(��z�id#"�r��$G�Jz[�U�Y�ǾQWO��]E�f���_�g�f�\������P_�4Y�Ȝ�m���#���,��z��ӂ���"�%%!A�B�����2��V���������C��Q�Zz��$�r�"�vC�ᐔ���Wt�eѢ���H���K����U���ʔH/�7Ȗ6�Q�v@%~X�7�!�x���ȅ��^+�^��������e B"����)t��UdQ�� $H�7���q�M�4�!��r�Dv���yM�&fO��N��&=%Y)��A5�����mO����VQP���U
Z�d�*2�P����]N�} ����{Z����׃ך���1�7�b�J|����^U�c�;.R�1(�`��3m��V@��GM0��4z)�ӒV�~��:��.iʫ��	#���W'��ʑ�!w8����}{����y������/�K]%�a��bZV	J��$�0�+w�ˊ���uN�w����t��L��i��J�#hq�m.��\E�s5%�`����� ��0pd4P�z1���π���؃��4���]�x���d֞���E=;	}S��g;�/�1R��珘���Av;��|}f�$�B�شT��m��@�t�r�-Ї2�6%g[���H9t�h1ѱG s�r��\¹����m#��m;��RaSs���!�x��hz���=��s�=)�u7����(D�]F��1�h��C'O�T��[l�V��`"�7�&�B��v�.��	E�YE��oy����x[hVe�B)g�6�%��w1�Xwb2�R��B�`��8�ͼ��T��MP�*Br��V5�)�"�3�d�dg�'��'c�B�0�����<�&6/[=�a��!���R���.m���g�vIvm�}Zw�ˊ�I�T�8�T
o�Wp:��Fq�5i�<������x<=*��t`%mkBo]&��3X]Ƃf�s�:�p�?Mt����L�pTh��ɋ��`ϼ����|fb��_��:�"u]�M��Fa@�� ��q:�;o����?q��B=qW�B|��b��ra[�����R��0Jy�u��6��nۮt35��n��Fnzk7���0�l�]���9�� ����n��ImVi�#�[M�(�M�������( 7/qp%�����s��	�#�H}�w�{����EL�e9��+�9�����H���y�k�u��ohhe����:'���̖6�U�۠�aIw�o�n��!1�E�5��}��/]׬���U+�h�6�:���N��1a��Ր{]�4�z��^gtֵ��ژHII�<:�a�<7*�(,�����t�.9ْtd�74gЅ�Pw�ߓڡ��WԠRX�r�
��=$K�Ms��s�t�_'�8���(�b
)���^�Z��+1g(��4��?0�`'�V�.�'�'C�ߕ�^\������zp�d�9�׏A���=�/vK}8��?���8����U���m����P.
�(��s�|25l�{����K�|��t���i��u%�@C"����!��}�O(�-@���fS��k9Λҁ���X���(�les����7ps%�qDa����T�n5����q-��o�x˲�Zh�]cwp�Ԙ/!�!_��ŀ��3��du,e˭͠�ʽ�Y���坙��A|�Q��������"��u�ydK����Ds�����6�9��k^��0���v\�X���f ��iUte8p���]��,���P��	WjȎ����'�hm�?`D�w!��W+X�3-�?�-:�
�NFW�d韉�+>���<�xd��P�ː��v�XF����5^x�Q`��H]m��������v��B^V!�5��AH)ޛ��<X�Z�h-�ۅ﭅�W��?ܽeW]�-
!�����[����8��%�;wk���w<���q�?��j�ڵkW�%s.�����,����Z4�����V�ˏd����,�_���0,=���J��`��wn`��r��t�.+s�\�����l��E��ɓGj�T��� ����]�[�GN����U}���Zv����sZ�೰|���_\��{4@ &���_Ϋ���wQ6���"�_ңa��	�2�-�#&�r�ݡ�n�ȳi�Ưa�w쉭�ᅖ�pTuwu�i��1g�b�X3�h|Q Kq'����������`Ă���f_��{S�%�z��R�n�D*�Z'�O����O�J��`Ƀ}���_��>��vS�W֋�ǀ�t��KJ��i>�����G�P6�)�B�1`1�R�kQ4�����@�gno���|��n�㍯d5��<�Kǥ�5g6��Z����*BMģC��umɍ��'�K��);+�����W�  8�&�+�7sr��tE)&�m5tLۧ�{1���uYq�t+ҽm�����FKZ�)5T"9Y��,��*d�U�Z>L<������ɔ�9�ی�nlr�?,�ۀ�9ؚ��Z$���RL%8�=����/_9��40�DFrl��ܟ	�2[,�����"0n��'b�z|��^R�ϧG�f�eF�����S����x�՜�	雱���t^^/>��O��]��{��|~��w��3Q�ӳO~g�wB�Kӎ�uĲ��w��N�����'4\O�3ն)3R��ꍮ�x��Ԍ�_�?ʐ��)�i=�Ln2.݈����
o��i'L�S51��\�#�9�ĵ�Uv0���
#��ha\�y�}?2�u�^-ɔ�p�˱ɪ�Di��-qn��Q���7#g�n%���
'��;����`��M-8\=��#��]�T�kqi�Wg~�,���.

E����;��)/�u/!��,Q�I�P�OQA��,�_Z�Y�AM�H y��KQة��T�<��{�8��k%,��U�ғ�I���c��b�O�Q��+��2�Qo6�lP�y���B��+�t�y�������_��y��ϼ�Xۛ)��M ��a��.߂�RC�rWڱ��@č؟Q�N.�R�G�g5�;��d��O�x��4LEd5��g�>Z�J�jGJ8c�C��Y��%x�;��8���h���=�ϳ��\��bl��ܻ�G��k0�,��_7E=@���m/��6�kӣZ.y��@��j��g`�	�����D���;�\Xw�H�_	M��E�L��qg�o8��>}��>�r�(L.(:���F��M��h��F�&��]����R�,��A,�܃���m���;��gx�>#*jl-M+����"����Zr��i���C(��@����� ��h�xX�o<+^�><�7�~����Ա�Z��3Q7�'�Hq�Xtr�-�#��D֍ z�����I�D;��,�&��K�o��9��6#�m�)$�Mk@�ӝ�k"���ǔ6�So6���A������I���jʒ�pD�.��?_�Dϗ)��?�����J�葷+0!b����\�NW�d�%�e��@�x3��8�jiJ���wB����H��'xbg!���&�Iz�BAÞd�^aZ��!��B��
)���k���$�,s���*��w	JFa�j�c��H��!3 n>z�1Q��O��=�%��PQ��-&h��]��s��1oncۻv+��hq���QS'i$}%�><�&m���ᓓ֧�6��u&`���ů���զ�N�C8� 6���9>�D=(��<HP�c��9]�ss�&ep�(\v�{9���xԈn�eX��P�e��<Kq4C��ľM���z?8u\�)~p���u��i�Z�L���w�	b�5�.Cg�o �d6"3�e9�@�1�=>�\/�8O�h��}�5���ae3/�Z��P����Y���4�3�a�]b̭��u���^p�|��
o]��򩸚!*EY/ʨ�2,�\���W�I��zN݃�7�#�#�\ ���A�p+���+x� �6����o��&J�\��b��XT�Y���womW���ӱ(s6�����'�w)c�z��>��n�v��G�n�5��ƃ��d޿$#ґ�7�G����߫�b��AK&Ѣ��)�Ên�'�{G��:|��mvZN���̺���Śm�LH!sP+���q5=JeV	��-R��I�[�k3v�3��ɩ�}c�ʿ{�e��UY�3��&��~�]ZA�xj�G�T_�Ԉm��-��ԑ���T����G�j�	���N.�b\OX�19^�M�Ψ.\�1��D�Q��1��� �����_�6I��ɗg���;V6g�0n� u�3�˺����g��g���5���#>	�<q6Ƚͽ�*@7c�'g�-�)ޑ��	�P��3/
�i=���OE�vm�"��<YEF״v����7��E���u�&�V]�7�����.��'ؼ�Ndm��.oPH`Q��z�f�3�������J�L0�#�/"{����j��E)����q�R���#��\�������aG-�1(|? q艗�83���Y=��J��nc?����}Kke�u"�"�=s n�m����]��8o5ϯi�=!�M7,Y"Kɮ�[1�.-�DM@�4	ٷ7�?V�Yoڊ)Ák.:��JNP�ʛ�]e�wǹ�*���b��j_�=�:�6�wxT=�߾����8�w�'>͘��0j����3^�=���?~�ˉ�濄<��҈��fת�������/�(P
������j��mu�X7�<��~y�݌�~��+eud���?��Ulܧ5>����ab�s�[�����Ű�-=s*Gp���(�����W:x�Ȥ��:�ȷ�����)�|%E���`N�溄F�A����p�n��u}��3�y�����?ܸ������Y9���Q�6��z���I&5`�����~]}�'9u�Y�b!�b�l���p�B  �1LrO.�J�`(�O�]~�c�T��NH*�?��b�'s�/r�C*��8b43��
X|�����Ri���?����`�v+(��a��dD����Я�ɱ��"�h�����e?l�5+�7�~��:�&~[�}���c?=�! �U׋��4{�V���[�J��8����2��J�s�~#�K'�ǶK5�S��yD�: Սik���N�")���BS(\)�`DP���� ��^�!v�J�F��L�Yw/6s_��W���d�v�������S�Vs�ě�����z���[��M���Ȯ��ZX����dh+����a��J8�EҼȝ�0���}�Y�<����c �l�0����J��S]���}x>��ŋ�Qq�ý�|6	��m�?���a}�jo�HbE	KM���d���)�)����A��𰨄�DW���-|�2��e�^���8�"���������u�-�W 	�Jl�֗�@�ЭE��S폴��԰�Dj���&��g��#��<G��p�'���QJzzD����-���T��0P,���{veǅ�B��w���,���`*ɴ�d�gR��D��""^�˷g,���ۿƬ��Y�?�&���X����N�櫪�f����Pb�\�H�m�����=���Mį�a@e��nk�L�}�8Wt�陙m�\tO��� ��}�rż�22������;ʿB�dB�_�v+�4�N�Y��Ztc�����8�J�R^p�֐52^���(l\Í�m��4@��a���<o�MC)7��t�P3QU)H��P�)o� �"�.٩�#/}J��U
��(75����X��Qk�{��|̍�Ua�ճ�1,���a�������o]r�6u�(�(���J����&��g�p������C�ܫ�p�٨���K?�6X�Xg�K���ކ{K��P'�:A�]*`�e^2�o��"?��y&7{������/%h��!���z�uO��6'}��|<�ќφ�dێ?U��r-o�T�T���{�tIO�'#��ΰ��JG�V�ҟ��$ ��6+s|*�i/�ź+�C*���	��cզ����s<���?[�p���¯Q������+>��g�(�%g������D�1��G�Cz���� �V;i��@��ص.�¾v�\���2H�g�!Q뚻6ߛ�]-3/�:K�t�֒�&۲��9EmPd0#�V}}M�� �Z1�&���&�Nn~�m��
c�
����`�t���G�R�����J!��O�7ZL)���$���k"}Q��l�[>5�$��F�����~k�L��bv��N�{v�@����2I�� e٤)�po�/t��6��&�]ӽ���EZR*R[p

���ڪ|�p�X��� ckt����@��}b>���D����� �m�CF9�bz0S&r�嵲Ϟ��G=>�,�� H�,!���`��YkJ�"G#�tP?ReǼ�����N`m'|�:?^�;�N� 6����a��ֲtn�@���׹3�0ux����c�-�7��K�f{6�]��tZ�z�6�a�yh)�j���
�r�M��41���i�̝G*��3-|����G�~::o��5��5� Au��_�?�z�I����z$���X�ބ;����k�w�������5��28���EC��V5{����},P��YOר9�c*���� ?�;,���{�b���|r�����1h�����Cw&k�Y�|}��!�5���r�1��>�֏u�{�L�G*���=B������nӦ��q� K6��ѝ������L��($d��GwY3I\�ګ��i\D>��ٝ����c�NW+��$�8��!Q�K��)�H��(�_a�.��������@�D�@���MI?�yE�c�l<o��s?�������l	S�W2m��7y��O5ao���[��4�YO�A��R��fj��T�Lz��^����]��lI��2�*�5��ơ�3���O�b�.Kt6����!5�=���nC��S�=[K+���GK�^)�a�0���K&e]ŦB�8gqTF���'ڊـ���~��9]�N�^�n���A�G�D>�.�(Ŭ���k�b�Rbd��k?���#��-6� ,���v]�'5��]5˕
Sgʁ};�+�)����lm�� �t��5~��a-��WέI�cՒ7���#�����1 ۖN*s��dg柮*�2��JH�-�B=�a�0�,������Ж#cclL�9��;+Bj�ُ��[T�X;I��7�93_3���кT��$≘�������F1x'E�\��a(��fa������3b���]8����7T��^�&'=τ^�,������Mc(i$7���1���}}*d���?��z�tc�n�V^s4�6_y�;:��e�nζ�]�����{[A3�؅�W�������x.*��FO��bb��"y��1�zN
��cƧýC��<|eo��7v3�W�"�7��B���(c�����#VǅMr$��=å�d������P����=R&��Whڙ�Ɲ���54�W~I��x�8��N[a|hE��H���|X �a�:��� O�Q��&<�l���(���A��Xx�Xۥ�h4�ӛ$��ο4[���>�~�.l���D?�V�*@��ȓR��G�U�&:����4�SQ��|	�l龑H��$b����ܦŎU�1�:]���D���}[�s 푸�z��Ց��ΜO̔��b���l���V��4�jY��J4��	6<)�HO�6�fiF�;�]��{�qD!����b�k���$��V<��#�@/(��Ry��Tw#���a�Y�<�/�͵��`���Rm��6�ɹne�hOC�32�z�*���~��\v4qd�N_�+)��.ϗ�+�n#x ���R�~�nl�ya�9h����Y;j�u����/0�Ð6"��m�5�e�% ��ju�K��`u[��E����ӚR�?�S�x@�ж�j�7E�î�[̴&8o�l��ğ�]d�q]W���\*���|#o�xULQi�z�b|�	&8�g�;R@<�*&�1d���#!���4��Y�f� }�d��V'o�'�3����p�$
��H�Q9]��܂{�/D5��3vnZ�����S~�Uu7l����ݥ<��=p�y����&d�6TX�]�U�a�Z5�kDǏ*�2H�ˆrT�X��_~RU��݆64�ĭFa��1bx���?oF~ra)�w�f�
��^��7��N>��p��ek1�IOΎ�[��W̤e���uP����n2�Q-�0�hI��C�|�B���w�u��SU�[i��M�sA	,�n���
��\=�xp���m�ez\�Q����������p·��2�"O,TPM�9��k|"w��T4<����g׉'6�Pw<�`�s��X��B=@��oa��_�J�
���M��*ٜ^hV��X�_�<�&��=@�h(�4UJ1�"%�W������l��(�6F�T�z�u���ul�-Ro�Q�Z4&�4��:m�GR�QT,��`+��_D���(�U�Ԉ.��|���׾0��nk�&�	�MG�w-r�b��{�P
�𓘫!�E��39xR�q�n�^��~���	p�ُ-y����B��jM����D�í2��ޡZ�?��c��I�
�2����H�C�#N~'��q+��é��ɑz�%e�-)��%�����?
�mMQq���+P+��Ƚ+!� 7l��ڪ�М�F�o2RP���;})dE˳����)��)	�M%%���n+UĆτ�[���d2V&���ZB�B1�Iب�V��]�H���Z�^�V� ����'^b�q��pH:�1���4�rY�"6����0NO9k]�Gh.#O{Pr��b
C�x�ф�	R�"��U�'k[Y�_��y��'��gz��?�֪"�.Qȹ���|pM�`J2gڴ��,���A���k�'eM��ڃ��¿�'4Ĭ�3��p������1��/w�zڌۃ��[���B�H�U��N��2�)�ΈR���Ř���&��]%���&�E�+�cܨ�T��,��=l�h�\E����O���a���o��M͜���Qȕgc!�ii��\D���m+�D��W� ���{x��k6T�/�n��/	VνЦ�}ƍ�K���8�_2�q�E�� ��F]D
k�h���A��L`��t����N"$�6�tG��r%�K%��h�U�gP�4CE��H]C%{x�_�)��{E�'8f���l�	i�twl~����O����Mi�M�7�'1����U	2v�}�q�`'s���\����Wu�������@����uB�a������S���������*��<n�:��QʨLӱW@a�0�e}�Wε�	��j���#���z}��Y>��d��Q)���E+B'�������5���W�4�N�������j4}� ߦ�X��3�eѹT�����"�e4K|GɑM^z�L���Ja��jڟ�
7 7�g�.�È�G���ޡ?<w�67�ہt��D�l�Y�ߥ�$�U�,2�v~���_w�#��g��t���uA��ߟ�L6��Y�Yu�N[?Ω~!6��)�u<�r���n\��<*�2����u
$%�=y��4����3�i��=����;�f<N���SO�L�����͌B%���Ƣ��|�p����I]_���k�	���jw���;k˒�'������>9�Q���-�7�<�G�0�w_�w��*�u2j�Ƈx4�c3!�����H�T�`*�������L�C/$��>�c�Hn_;`��?�@s<�1a$r�L��UU���uF>W7����;;��p����t�\�,���-�u�'�zU�����k����y�/K6�Eμ~0�Uw�dnmܚ�4����IR!�������/���@RC����L��3-&w ����G�L�V������p�Mޯ��Oe2�dg�`�Ϻz�v q�[��|��U?�u���������Ǝ�oZqh)qY1�.��p}O����  �;3�ŏ$=��;9eC�=zw�YU��ԔbD����]�;^zt�p��%�˹A�mo�H���r�y��6���v���o�{��)nX�y���o��&G$�&�<��o���S� �@��0p��m��Q�K�	h�f���{8���2�I�������W#�E#�A[���$V�1��A���`�
;��`�BDU?ۦc��C�*jO=ʬ/��x��������T!�q���L��N�G��s"yB둻&�Z�e94.0k���Is0�쉏�:RGˑ++��@��Tp��(dR����� ��C�|���EA��_޹C����T?T�Q�a�}O�h|E:Z?���J)#��,��i��'2����2��;�ˣ�_������f�0_�.BfQL������[`k0Z��Ͻ��N=�J���;��B���'��W���ݽ��ҥP>j�rX��=t��Ü�[��H��J^�n/�c��K87�|�<,����S�C��7� J�r��|%��S -�HD��r�
l �$�/����qײ���ޘiP`��ԋ��xk���YjWԣd���c�ݗ��_'��\��O��������N�r��O�9�=�%�~���]�I��X�_�`��%�ߦ?�'�_Φu�y����n�󩚒�q0�`�%k�cņc̋y8��]���μ�/��P�!3�\�u�C�ydol,��B��Z�C8�du;�[;Ox�|�9����<���M�[�<N��8�Ɉ
��NZ�͞��WX(�EZl���e�� j��q��S����#7��[ackwR�)��ɉ�⤺�R̋�<p���:6;���]JS8l�`3����]�-.*Ä�2~L��~vW�l��
WQ�D+�jO��F�ޜP���j���b�E���6�!k�j�am�Q�GLX&A&��Nk6k����R<�I�},�R�֏m��Z�8`ڐ��)Lθ�??���p����n�Ӂ/<<| A?G@Z˅P�~
n"/�(�e����5`CEn�!��
\ֻ�w���Sm���
�Ԝi�J��������2	��W�%J�ox!a�%���"�����J����d~�D������yv��L��"�2G%�{Ώ(����I/�� Tjo�v��{05w�G���Ų�?0'�(M�Q�Yg����h�;B�z�U)<'�g�����fh}�l��	BI�Q��ٱZ�vG�����ez�7<I��eJh�(��̂��۪߫���u�sk���0Lʈ��0�"��H)<a�A� �j��妫.����>�X懶�ctN'�xFw�+}�F3b]�v���˵�������*Y�D�5ԏx�kJޞ�}���^���"����<��'K��Dm�_��|X�۶��&u0�F��销FP�����`S�����&��)2U�o�]���]�2���Z/�	,-���,}	�����ή�]�D^'~�bŹ�V^XAG��K��H�Gb�/�)&�q|܆| �'ߵ�QZ� Ќ�@��ɵKG�F=��ʈr�������e�n=!g�5|�-d?_F�(#�=�f$-;��S�U�-�mk5}d��;=33��~X���9^�g����` �>��~�\���>;m39��������~Ɉ�2B�'�S��n�م"{ӹ��l+���\��=-���sl��!/��3�}���i�?+�#�s�q�n����+[�}��4����~7t}�"� ��o�۳D�鈲m뜷��Pw�c軕�U_��h
�����7eg��#��֠#���A�(B\M�E�z�%??��d��xc<9lΐ�Y����V0Q��;#�.��a��Ą�T���9#F�d;k���-���qx- #��3c��Յ�ݕ��pgn�>����)A�V���N���h�na��*�Y�sz�(�l]2��k(p�
���� .?d��Ҿ�N-��8�ɨ	�F�i����c�1��)4{1�S��b���S�"�KNuy��x�%��Zg�;n�2Wj���{h���ou1�s�B�^~U��\�\v,U�.Bakf�0F+���X]�/|�y�� ��% ��@���'b+�ք�d���{�&���%�(ڭ���M��q���;���k
x����*+��:tY��Z'�3���KAp��:��y>��f����1媬�dQ�%��Ţ�L鈘2�a�
ݷf}RuV�)z���/���EX����]�x�VGMR���I��ӂ�ŋ�T�>l�(8ld�w�a�5`�?����Wy^'�VW�Dk7��d�6oX�Lb�9�U;Vi�e���1���#F��nו�6�뿅8F:^6|DՐ�O�)+�>>>N#��(����S�N�͓=%�����n�rP��O�,&s�}�|�zX�+Ǯ������'K�&vM�k�U�D�,��g�_f��^*ړ�f\ppE�L�^�u�e> ��v[2����&��� ���j�,<)w�k��d֥�����7�Ӧ���ʉ'�zv����v���4ut�U^V]y����uUbMw3��]�1�o��߳�۵�Owv���ςܷ�����j���'�k�b�� �:W,�̉P�6I�eֶ:X��\�mjz�q���oKPi�����C�K/#R�Q`�P�(�,�3����ta�`>�3�d�c��P�\JPwi'�d1>����[^��߫�"��3��F�~���#���_�cR艡N9P���4j�}�?#�W���12�/�A3��Mo�e�_����\�7l����jl��re������NXfd�"��>�zcJ����@S۬�.Y:r�c�1��d�OX��ti-;���@q��Ϧ>�鋬Ei��z/?Lfp"x�F��_���7��C!	�нp��)��!�֙L=e�O�wS%%%2!�IcWX�Uݨ�g�����?!Kg�<s# 43�1[!�A�mԖ�o�F�m4%
v!�3����G��C�+u�����!�U^;$�C9Zl�Q�[�r@hB<E�Uw偪n��
�*�Z��F��\\V��M�%s�2e5/%&�LT���A˸I��n��TI;� �,/3$���]=�skJ���a�Z����8�ߑ�4�-J��%�BT�%CQjCB�|��g{cx��Hl��c<	ӌHvT���F������O)&Y�/c�υ���af󀤿��=����W����ɋ*X4uy�Xj����D�Ogܷ��{��7���CM�N\��I	��e Ϝ�A�hO[p�P��ڿ�T	r��堋�	ܻ�<b�=�/$��- �H:�����ݍ��T��$���F�;ل�~�%돲i��E�?|�nh��o������7��uT�zq�$n�h��@���H�E[��]���ft���ag�����c�&��%��t{�n_��gܒ���2mْ�x:��#FG�(��=�����|	� ������${	y[���!�Jd�>��S�Ѝ��W�Ǘ�'�V����ޟ�P��8'(���#����4p����h�b�h𝖨����}�+j�ϙ����t�����K���u}�g����59qW�Y��Lj����d��_�Eo�Ǳ���ֵ��n�OK{7��A�j�+�^�ࡘ�Ԃ���QV�Ek@��:=�u���;2*	�]m���H�P=�i~Ɔ���* ,X�D����Ҵŝ{b�JJ�����(��G����r��6��̙�sq�T�3�R�e绩)�j����\��7���Kag�3�q����\��8�\n�dc�f�NH[�S&�!>����B帹����8b�����@�)�<�VYL���)N�{�H�T�SN ��ty����Q�ҩ���M
�ThEe!{I(���_�r�a�⇇�_�fwQ�bq.S"��w�K6�"E���~��]��b1%�-
hqM8��tĶ����W�Pl�4\��-_?Vi���)͵��5���;}Ж��2rv�kKk<����j�$f��E�dT�R#s�(���V=�^�t,ǧB�b�ۜY_OFZ��n�Ӽ+q���B��Ƕ3엙�2�w�С�[}D���O!�«zIBÎjvl��F8Z+х�����EosTO�G+�xGR��h�D�bАz�?�DgvI!�	��Ӈ��OhѤ���f���kg��"���`Ǜ!��h�Di���d�,�N �X��:5Z���_�X<E��y�Nۦ���������R.Q���UZ(%9��p�^��щ��Yþ�P2�[��=v�Pӿ�����k��ͅUg��j�KnW@�Uu�⒟nU����}�Y���<��]�J��9�a���9�V�ޕ���~,_Q�bRpN�_	9v��������}��2}י��Yj΍��H�>�&b!]`��'h��@�'l.PAe����[*�D��[�Ǉwps�\{*b��0X�Q}��7]m�F&�t'��m��i�2�ֲ��[�l��;i���HS��FD��/>�/I�cҫuޘIn.��,��M+�m*Q7Y�x������E(�L(3������̘<��`���Uړ7.!�~����ƙn���i�y-��52���+r�
�fB*U�djrܳ�PrR���;��ø�:�c���C@E�
d�������a���J,����=��T�f�ˍ;/���k1���
Ӣ���3,�����Z���ND6������aZ��CfEJ�?{I�s���m���#cx#����yJ��b���=�^f��͋�������`�ɳ�_��?��ޝǔ&�
��˝ۯ�"�t(<!xB?�no�a9�t�J},F�8w�3�"�ş&�w1�����;��q���xt���=$��|΢���})��2�<�55�������(��ЛWK(�>����%ѫ�y�'�9�L�I��'�a�~��SU������M��x���z��Q�g��.D"Z��#+�4���]@�&�,'�h�.i�Y�_9�$�͇�i��ͼEݣ�u�ε0H�����S�n���M�\�+Њ�b{�D?T�~_I���<����]*�mO�X��滎~yz,�t8ð���e$p`�k�	x���O\N� �[\69���}��S�b�t`ēi�޺��������fš��L��\[5-� I6���*��]$����o4V@
U�F��*H�Tz%B�N�uL��my�g0��}�n�k9�t~[��f�kb0H��x�5�:�n��
̇�j����3�

���Rh��l�oF��4�0��u"���w�Jn3�wE�a�B=��7�����`�%]�	�>����D��q��YC �¿��(kQZ�O���2�mwx�O3�ʉ��X.�t�"�����>���y�!l�������G�L~v��c�A�˨�B���ƖyI�Vsz���A�m�ū����]������$��
��I�=KiE�U�m/j_�3.v#��(싆�4��r>^6zQ���(�Gpఠ�>��\3����p��K��~3�i�[u�H�Q�.�	�o�I�����Uku ��
�T�`9�P��:�n�B.qO̡���`�`�Ui���ԃl���<�0�i}�c[��A�3k`ap�]����O�q��t�����?�f�걩+�Hq���%}\���X�����x��
 �I���!�8�E��NH�(���|2���{�|��Ҳ���b:C�l���vt�%"��!'�[*��c��ޱ��S��`�wg�y�'Z��O�5mS�-�LVݣ����j<���k��$2�yCxm9P~P�\�8�)�+e��{B9(x��c~+��汯s�_g��˄���1J��A���CQ�!�_������}�㒛��s�d��~;P{�(��[d��`FC��λ�������	^�Zq�|��q��*�5o��_2���&��6�wQ�kk����ڥ:H9å�+�9�ׯ�j��8����E��U7��c�_�BeaO��������<�@��r^?��|,��Ը=<"<=|������O��O���՝�����-�Q),�¾��1�*��F�9�+�#�r򒑤<��S��l��X�󺍁©����n�S��F��K��⼱�v;�!�F��{��>�=�;��6���=���V�NL������Ȃ��%sF�����'%h%��.���Q��	�zt�T�����}�H�%���JIi]��t��_L��bPn����{8����Nhm�0�P�%'����j�H,�$:�`�E�L'jͣ��QYb�5:��1�J�ɨ!r�/���v�E�6�E*�����;��pS�Gh��,l�L�$�9�:�~��F���l`3��@�Y��2�6�.�f�$������-\A��ȥu9�Hs�򀬲`����J3�����D���7�&�a"�,�j��
� ����맪4��Vf���J�$��}�	�OzfU�F!SI��j���ף6��􂱴.Sof�NS���j�����}���9Vv�4X`�Qh�8v_t��hy�J�B�����p�mohak�>�fz#��n�����<��:�7� e��i�Վq]��X�9�z$X�36%����r�G������˩��q�$�Sf��)�.��F�ө��4|x��6�^R���E�a�6[��X��8���Sx�w��h�s ��:��H����[5��Q��4�^��!�k;��v���J�C�������~����#P��\��#<���vc�\j�.[Zu���l��2�ׇP��S?U?�o���ܷ��ޟKnƖ�m�r=�ȔM�~���ֳ�+��>�ܭ�� ڵ)�C$C��fc�:����g-����/d�If��NB%�zHfrC�7f-��hW��Bb2//��kGC��9)�Pd��/�\�dS�*���v�*r�}��Mq��zX����ě!pv}V��ཟ. Vs���ѽ�B�h�(��씎�a%o/�L�R @M�q`}��k�ZU��=9;P�/o�+����fR��\�4�D�g��|@#�|� E\�OpIf��Jj����d'Ľ�7p	4�����XW��ƽ�J	I���^pH�7��:b�b6���s{G�UoFGG B�v�s�!�sn����������L�4�K��5�Ob����5qa�s���2����'(��*挖4�q���u��ڻ�_x꼖F��D1}��a˱��)�KA�����8��i_�S� 敚E:�,�γ��n½`�fAw�����찧���#x��3����"T�ڴ�L�+�|Qo�)͞��7&��Q�%��~6�GlرFO<��<:
`�:T�����x�=+߹�vQ���z��V�T g��;�\�:[��@���Jz�n�}O�&���dV��>o�����Bk8�_�Il�ۘ#�/n ����wVd�͑�֯�����M�)�
�9�=c�k��4`���A'����jڄl��W[7�\������f�	�PwΈ�@���T>-O��x�奚�C/��3Z4����e)Z"��ByR�h��<���&��?je����Ye�n�*φ�j=)"�`��>�I��0i�M��%R��b܉�,MC��e2Vw]�K��;�kNN�ղ���?�B���yH�[�L�f����&�=:��!!(0�T�����^>u~�|��0IG��_����(D�8�ֿ��n�͙6��c��!x�2�"���Z/�a!�yh
���}
�΂c�:J����J$J(ϱ�V�v�d9��I��[��,d�?��1��/��-\�ϭ_�'�X�M���|E��_MyDʂ�� )�i�̙����#(��R���ֿ���+�����2����V�m�#RF�fU�l�ń7�@n5!փF5�UAe���#�&�#��&ۦ��Q{��0���&(�ݿ�(�)X*����W���NR����y�e�Qڔ�Mp�o*�]���pio�ۓ��~wK�."�z�9����EZ��a����F� @�D�R-����O�O}���N��]	8��H�Q��h�9<O�զ��0[=�yU��tx�*i�B�!�b�%!��W�&�"�72���T!o�0��3��]0�X&�b���G���  Blr�tEE5��
�p�D��	�*L��U䛰�%Q��=�]y�?�t�Z��zz�(�C$���t�.x��'�ίɈڦ���ֹ����G��'u����7KF��D<��)��'5��a��8HU�S�!��(�dx���n.%��q��)፞�ɤ��
Wܷŷ��1)��i˵6�9�_w��������*�BA��/���DC/b��`�#nY��M��ꏚw/�n�b�e����r���Y�����,?�J,	�߼Y���:T ��3#�z�
���EM���3�piDx���5<�(dx�;�"T0��H�3�A�q�}
�#Z����������pQ,��*ܽ�e�I�o����ʨ��`�����;'�3Xpw���m��w����%8��m�7��k���u8�S]��z���i�[>�+CQ '������� c�w�FF�$P"1�?W���$.����`b*��ю�a1���v�?0$g�J���a���1m�إ�0��Q�IP/
h�s���{aBd�K�W5̓7�n+U�%6�W�F�CgM�#v���'�w^��@��"8�P�h�g#hxAu��^JFw���Gj�Z�:�!F
��I^��[(�����	���Iˍ�Z��0�nzi��t\���vrJ]�!x��cP�^��/����з3S>J�8�(�Y�����2k���#'�n0g(�J��[a��։窗�^c���u�����'=_b; �LB���\��c
k�Y�kg�~�q�5��(�ŧY�����8�
_��Vsl�پ��뮥��ǫ=�/�FY�ղ�˲��}�@�|����^ۼ�f%! ��^y���Cņ(����I��b��FC����XBm�l�@k�?�A4��c}_5q�� ge�+ ��-f�&��:l&�|g�87
��'��Y?�m�Կ��>t$j�����-���,���`�5��k�e� -�>>P�>J���ڳ�S��We�,��+eg�������_��<����T��D��OhpzD����U�X�Z�z�j��f� ��/����r�X4n}��H�8k��MV�yzV�ð�TI=���x[����&�̕�����]�.2�b:��<��Az��>�]�ͯW8���=^�Gj�ϫ�tq�$B������6փ��H�	@��N>�u�G�`)�>��p[P�&�Zʆ�/e�~\���q2�����j5J��ˑ�/Sz�.\@MӢ�k�)+�Ҥ�e���.�a�*��|����t��o�2��q'����KWr*��݉T^�u�
��@}թEI��#���<������T��]��v?U�+�֜�Q�D:+�w,�21���U�V%2��X5j--�Y���ҍ#�Dve��������������	����f{2f�S�.[�{X7Z�h7���7:�$���`��Ch/���Qߍ��t��s�=�.0Y�[ P����Ks:���G<�Y��s������ b�o5�0����Ep��݅������ J�D[��<�O=�=�|�5Y1�'�_�����0Tg�M6 [�Y0�]����tW>}x��Y��������l�і��Vˋ��I�>s>vV/�D�wG�/Uݧ�A˓֒��˓2m	�y�\��K��5�4��H	.����;����D+���sf���4UEV�y�#�O d�:�l�n#8�d�<�W�!��4�P�D��m96i����
��|�@��?�����I�����|�ח����dK^����5��P���kn������4�֓��#B���s,�z��P!0�N���3��q���L�=v*\Y���}�w���=JnwqÆ}�h��,��.d��zE�\|Ӆir3��|���de� -��'9���	XSӽ^�&���ŹmU.�@A?�����ϟ���^]��vË��6�mv
C�O�OA"���[~K+.�T~��̍�����\ �YX�R�p��8�}��@P�]
�b����
ٟ�__~ɼ\*t'��1�m�Ęȟzlo��_a�
6���G�-�6�$��}0�ܩZ�.I:�{���؄��c��F���N�M�G*f'E�`�Pi&�dM�<bLV����h�?8������!,��]g�N�%wI�1A_t�1�����*W�\�My���P>��W^�m��71[��@��Vӝp9�z�Çhژ�}瘃�QvC��^���4��]]<�c��s�5����������m��z8�{#����|�Y`�e������ /���ib���t}�cBN��+��t�S�ÊJ���_8��R�F<0Ҳ���B0�XJ$Z��>���w~�\�F��>54|��9�U�pZ�;{�5,��H"SQm�w@)�UT��������߫��7"�+�7;�c|哘4-�f�� �3 ����^i�j�I�^���Jx��S�x�v���A��V���:�*�ز���C1�芵����U��\f!kmF�_)���W�e��d�S���n�ݭI����|~���0{$�^�
��`���ʹt�7���}3��c���U���OM�oP���������������mt�z�����]�Z���~up\�.J��4*YϘT_�Bv@)��x~к�̃�S�E�w���Ц̓^EL�!���UC���bn^r�w��ʚ�{���2����=;��n7��O����܆m���Ɍ�O�*�©�ێv.�m�q6���3S�E~)�Y3�%m��n��U�߼���D��|[����٣�׏(eg	�t���Nbe�<�J�d�ߵ;�x!_]�]XfHZ�`���&�dBLh P8S˪N;|�6��tG�Q�-��y���jǮ߫V�����$I6���h����(��~Y%e���T7r�@��|V�0(�ų���V���]����	��J���/c���)��Z�Dv��(d�w�{�Rǃ������F<NN��Fn�u��
S�ڇf�w�%gs3;��(�U]E[�Xa�� >��Ou��cLFȣl�:�DC���(J��W��ɅQm�̀k�dQݻ���Av�W\eJ%�_�)1Bf�:�����j6s��i�G����Pr�&u	f"˷1Ҧ��`�Rks�U�Q��h~x�m�4�0bjg�]�Ql��l>p�#�d�%/�G~�{��ʢ��崢z�H+6ߙ�����.|���<Q-?�:���2���x j	��1}�h����5+I�8�$n�~w6�{.|Z��s�Y˿V�+�%|m�E��2��[���dq���D����fL��,�l�R˅��S��#�׃W@��m>��h"Y�$��P�� �E$���ov��X���N��42u�u5'y+q	�g�K	�B���b/��͡��A,4��BT�iA���x��!ֻ���$f^ޟ?�7�$2*[�.�Lz����q#���Q�t+v?�C�b1�z�����(�q;�A/���	�n�2�晴A������k8��H���y�l��.�΍ů3��t�*Px뉖A�D�.{^=����G�A%Q��#1��ϸunp�KbQ���N�㽍����̉?���T�3F��i0���	fO7V�Tv�s�w=�f&������c7�틯�`Xz�d���%Z��yAP����WJ��+N�` h���{�t��n�3�X�]����Z�Sҡ.[��B~���i�K��TӍ8�x��yO��hL�j��}-�����A�e�������wz��5�UL>_�ΙGx��zq�yM�4�ɿ��91�?(�NZ���_|�k�K�$V`|T�S����a�x�C�t����q&qi-@\�fݺ$#�����<��}w�(�y&|�
6�5=5�w�7�]^+�|f���{g�n����Z�4�8�l�e������#�ōbP�3�CI�"O|Ż��A�VG[��;ߒ��C��`�j����!��k�>Y�s-��.�.sc��/��R�#dlZ���3�w���ߴ3ւ}�]<�
ġ�]ᔍ)������CE����8�<Z�/C��,��B���^���-�ҋ�j�qy�pOd���k��:3\��"J�t����t�X�u+�r��P��<�Q���S_��%�pV�e#�G^Ek�8(�_���%.�7����t\�{O�'=z�����j��L�}��Z�n�9DV5e7$��CJES0r2�T|'n͚Zs�^�����Ħ�	=�	W��e�����.:�{���L����Ra���=i�Ǩ}�A^-�HC�S�@�5�AG�g�[˺ν�D���m_����=+�i�۟�\�an�/�b`��1�L��%>Jݕ�*�Tj<�j��_�SP�G2yu���7_�*x�c�H���>���Ӭ���	�Vu+��D ���n)$��4D1o�sw)�7��ҹ�$&��/�|��E�hyX�IG	�FFe۹M=*���s�@�d�뾘���%H�n�?�T�p�^=mn���I�.��<d\��<,��&��>.ΒB���_�Q{�<4�l�X�t���;�|?�7���#+#G̫5�N���(�&��%��g���ٷA$H�>�
!缁�1zZgFْ�. �	�R'�B�k��8̹�#����V�4i�����(�O�2����5��C�U^�8��
��G�����h�yJ]-�#��bJ��F���nL�
��N��Vv�MF��p&�M�(J�h`�1-�q*���#`�����<�6缭/
�T���F��Gb� ��&��9^�3z�g��G��&m'>���L�V�Ӝ�i���K����K�A?	����9y[.[��u�f$
�W�3�|9�<$NaIK��$��T�<rד�'��,���3^�'n�y���J�Z��ld1_�E�j�5���܁�=��K?��4! �xH���<a�Z�wBs^�=���QB�Z��1I���f�zo�U�Vw7*����gjԐ��ʆ�s��T�\?=�C!��8��Ї�
���8�������[N$�(��F$B�UQ��c�w��'�e>÷K�����œRM; ��O���-���Oz۹͵Zթ�:���#��en*�EZ�����ļ�.���� ��	����K 'e��ƶ�̘���צ��ء�S��$�D#�e�{��<�R �@�7�ޑ2V�t�]M������/=",���.�_{����4��w�����驕sn����j��ڽ2iPy�ė�=�Ϸk���$Pu�CT.�!H<�����^hB$I��r�Yt�xl8[��3s��od����X58��|���<g�R�;��X�
�)m�� `;�ܽ��-��lT_��E�1��q^�܇̳y�2C�`�08���x�[�% x��矉н�D`�\E !��lJ�k��� E�5�Kګ��6r�H_���o�:J.#���e˞�p�<>N��Q�Gb�ɐz�:�>�)ĺ�I���b���◮�u7x�H2n�Un-$���Wi�	p{�0���_W��y��b>��.�8_��}WD�f�����<��.0���U3
,{��X�=�?�E�u7M��J)�ZÎ�Tׂw����]p�C�Hd���S�g�kcu�@�u�
�ǘܨ�DXy_�#�"����#"b�q��A��vq^���շ$c<zo��VqT5���wm?�+�����N�.�>b_�����B�$��h=t;漺pu�(&����o���s�u׹}��HG���Y��G�P�/�s�I*�,��Z>%��p�@���;��qk,1M�N4W��:8~�iB�0��@�����/�/���������5GOh�|
�k���:� 6�͑�{b*k�ν�,໶��s~��^�3D����2�`R/*�A/Z�?9F*��*��*}l�ҭ�5�����}���W�G4�vE&RÝev�IJF��?��@��ǁ�Js)�g��� ��­�������2�155�_^����NMb�S|MՀ�{O��M���W{��k8�ɠ����n����l��;�n,��3޾�1�
��;T�����wt�(�n�ʎt��O���H��h'|0#9wD����f�� ڏ�/Vv<�����Y��ާ��W�*�2��'��^&�)���Jx�=���N��4���x��IZ���]��>��;,+�7�2jeD�`(��07���G�MTt-�M��#���ׇ�;�H�f�c�4z`���tI�����v��#n�I_��/��K`��~�s��d'�\��AP����b���j*y�鷀���n�4�R����$��\��
]��^�2ݬ���{Օ�؟�0JfN<�����C��f�	)�k�ɢ��x�� �����[��,Q�)�p�h����')j�;�l��31=07K�5O\�\���-�	��%YI)�M���l����z'���l�s� t�MMX�v�̐�<a���L)����]i@8-x�ZA:"��JX N�d�����!o���`l��b���X��_K�Ą2@�g��/���A��+�XYB~>*���8���;�b�?KҵLZ�q���?�	��ꮶ�W,�J�%�d���4KO_N���)��.fՋI$����n� JՕ��0T�d�;��W����n�Q��e�7��ŚHw��H��O�7؇)���ꏰ�jw�ۘ��ӡ�>L�nsQ"�FA�Ê�����$��9l҂��NaB�0�= $2�с�<���p){'���J��(fnm�������d�5}�e�|�~��Bd�xb��6��ѥ���R�
��̘�^�W�a��W��/����]��.DB0X��� ������H�I��N�Ő�@^�]p�Lfx�=J3�C��+�NS"`ߩ���R���T�rȳ��0/�/��DJH�_�U=��$ G�̹����?X���D$�l_�r�@e��`��j�Ji<�	i�UluHI��|��%�t
�Lݖ�J� ~;"���e��"KLN��'��CTu�u|	�o���pd'l}���8�|��� �7�ܿX8���
C \���fu^"����+ �X�!�ݩw��ey����B ^��Wp-g�6��[�ȟ__db(�r����m��::h���:�n�<�vxĜ-����e|���L�E{+X�۞Ɍ��3���J*��b�Ƭ^��I��5�~�&�K�ss��I?7;ҊP������+�լ��p�0\0�3kz����?��g�Zx���F����g9�+�͇V�DP��q"�k�g�d�t���@�P_h���P�e�#�(kL����2zذ���Ը�����|<��3�1�tf�$�78��󼨷���J*��0����e!����l�K+�JɱɃÓ���'��[��/V��������!��[x@�xX$��O����Q��ݼ{��Б�K-�^�u��dd¨��Դ[�h�+���j�o#���0�D4D���SvG��ؽ!�1?Fw���
kڥk�p��I[�'a����O�W�1�Ę^�s
�΢6�\s��hr�3��΃N��
��͓v�VA��-�@���Q˳�&.wGt��P��U@�;Ǩ�1����ŝoq�H;SՖة��n�j����w��Jm�@��~D�O���>���_H0����}�Vv�5�0����L�	6bF*�L]8M�+#�T��u4��8_��A�!b/�u]����@�6�@�����-�1��d3��]E�T���b�d�C�_���;�>*���t����\z٣���,d���j�f��@c���B�|������RK��@�oP�`R���`�ʰb�����<+H��e�P[���*��f��%{18�M�V7B�Чx\֤y�Q��ZZ.�;�ԌRB�F��w�U�$�0��AZ���.���,|9�B�|��� �ҜI����J�ё,k�?�	䶁������վXN���nհyI��������4/����JA��.�&��z��~]�$����� �E�_�H^pϙ�e��^��䷾p��Q��1��\ �p���$:�m2xa�0t�&�K�1�X� S��'Vo�"�L7!��t�Ie��q��V�}��u�Z��ѵ���o�`M�S�U��@��r�(�����@�)	 ���|����ߠCm]�<�>x�U��)�\I�3	��Yi�wTྏ�<�Xìqq�t�+�����yL����Z�����F�R32T��+��>��!�R8�o�y���Y#�G"J�Y���^�B?4S��mmQ�݁4��}ZtC���S0CH��f�F�[Ưx�+�"��i��wcO$��\��.���iwj�2�M\����yi�Y˩D_�9w.ʱŎ�
Г��yL�e�(d�6���@���2���-���e,��?�������#��F�3.�Y���S�<UI� ������/�;�������n�<�~( �w�u�GW�{�i�����%�c^%a�m_eг�<)f�q�R N�J���*�_��0��fp^�S����U��� U���Z�D���JH���EQ�����j�Y����c5�����5�D�*_3��y׷a��#��?���״bn�bH%7���B�ʄ�u�}<H�4ij5}ͻ��@m��`h�e�@��q ۸�]ٿ��0lB�E�Az9"/�;�7�ݚ���� �<.�s�%�^������KZ߄U�PRv�_�ۼKU���Gʇܲ�3�j�Թu'c�'���-Ӑ�,�ߩ��L�l�	��m)�[�\�`��y���,�I.�T6�/���uU�@;tC?�en?C�[��9P�@n�+��ő��,��������SP5����W�uv��&���d��Z�B�缌̱�c�Z)l��1ãz�J6k���t��	�����/"�	���͹�j+�8y�s]#�k��.oz��g��!��g/�eп��4F�rmxz�V�K!�{{ghMǇ̙���ӎ�Q��b��2I����4�䅘6�@Ե'z�sT�Z=�[@���>��I��	��c~��8#܂����/v��b$�s�6LG�"���z;<'f9�Y"ե��P�\���ӻ'��8�m�:P�>�������о��ι�Zv��i���V� E�dKr���x4��X�4,���,_\F�L젠��X��n�Q*$������x��`�.�?��tV�-�n:@G�1v�|�����|D��7o�$/o����$E�+w�=��n�v
������.'30.�50;ND�}�O�7����'Fj�>nb��Jh3��� ��"�D��)�	ҿ���Y�啧������:#!/Q��~��g���0�5Y�39H~��W,Hf�*ȝ����9P�͊!�MM9'� ܃�8�?_�o���6.9�XrN�Z55�Ʒ	7U,Vz%�d:��x�M�mRw�w�k++��f;^!ưhuVR�8��|�d�FY�`#|����!��������9��f�~q����nͻy�T�o�B!W�u2�e���꒐	p �翐�J���_1o%�9h��"	b��zs+��;OJy�^D�%8s?t��Q<�}�J�h�bp��Z��(��[�b��������Ɗ=�xºG���˃��)Nz���U�_��ߵ��Z�۲)��/��DL����Α��>wkW�55s�./L�~Α\ϣ�X�ƞ�;t��!���CB$��J�|�|�٥L$�(Hj�/���~�.�K�B��Zp����|RT�� {j�"��Z��H"���d,�Vu?b�ϔS�\zUB�U?�ɦ'���s_�x6��zw�H�v-ށ$n�ކ���J؃�fKO���Jt�r��n���U�i�����r��JҖ��>"��47�^�U��q�~��d�{�Ó�K���:�����ȋY�7̐�ſ�G�h��G<��8�3��ʻ=��롪fGFN���W��h���z�p)2�Ϟ��_~�w[<Y/7���#~!úU��k:�I�8��n^1Դ/8~�a�z� �;�{(�8����.�$����#w�4;��w�����"8�E�䗮k�Z�0_�l��s���_0�TA��@>oQt.�ΐER�r�5�Բ�®ܴ�Oۻ�3��-ܴ�4�W�?&�8��qW������,�o<�O�	zG��5��������m��~^��3������^�>l�F1/
�|���\c�$TC�i�ß�2�t��ߎ��b_xE~��5x�t�R�ة��W\�l0.a{�ԝ�w����Y<��#��cʿ��+$.	]b��.G�^>j1(�K	�����	��rm?T���ZjCaau���� Q}�c�� 1�����l�Y,� �����r��M������K�T.�g,T"��тIzv����<����;��ϸsng���o��w�#2��0�Ǒ c���,����܉׵��sLQ��^�aK��뻟��
��U�k+9������*�q'U�[�&�>���jml�W���Iv��E
J]{��S��Vj� d�0_��J�ѥ�\����_fs����mWE@��Å9K��/7��I�%�sԫT$��Ex���rHgFI�b4�s<�$�����?'��>������ݘGϷL&��o*PS]�����G<]l�DS4�����(�J�6?]V�Z�Dl*w��OW��ξ�x�vŕ#���(w>�_�p?|��{\<�	���@"���q5�5!�|�v~�EY�XE�|�.GG�!��^��i/�mP�Q��8m��^��n=O�)���x.5,����D���z/2l�r$�����}៊��:������gE�~TcM�_�oFm�=~�	�D
�G�^�7	�/J6��;��� 0��
��S�<�r4*h)�gc�H�B��|���lU%�����=rT  ֨"����.��d 4���[�H��1�4�TM�J(�իzArp
�wp��yNo���M6�]Y�&��b�k.E�)�hFs�%_�D�6���uE����Q���\�����+Z����)t%T�mX����tb:Y9�;b�>$Aч����U֮8����Mu�m4j�@Z�K>��.�O͙������' �%��?�˽�/zo�s�? �F�T�.ʃQC�T	�֫�ڭ�g��fA����K�2W��u���)�4�M]K�[bD�ۓ����!�L�/�]�u������ӈG�RT��������w�n��(�HM�/���*��a���&��7L����0�A	��a)Dگ�:����ЕD7e��n����6.�0�6�
���{�Ol�7���d��@��L-�:H�<<��+�
nʷ����1w��2�N73��\��ZJ��6���;��+��r���b�=�	i��g�8��������-��g�
p��UW#e7����vR��- ��%�N��|��L5�/l��3��t4��U�](�?�<�{�h\�{�|����f��9��T|Mb<yj�O�㾤�b�0._��kِxc�J�K���|H�����2���*�&s��IO�"��?k"���1��٭��䈵�yV���M&|�!��SB�j���_��IoHp�dg�ڿ�����
��jy=��n�T?GE��G�D��Y0N?,z���Q֓��{�&0^{9����,*�_30�A�h�^�h��R�J|p{ot�����{B��?BlrXm'f�]'���]�Ŧ�b0�$�G���U�[��׃��x���:�fB�W_�6u��[7$d��\7<��`'y\�#�_���-9{SG㈒
�:���ln���U�������>����
�@Xȍ�G�_��
�?�IE>B��f2fe�K�un_P:H�V�HW�ى��Gv�+X�H�:a]Ye��5�̥D�ivq���%�����CCAi^�:�����oA����G�g;6/���z�%��e�Z������ç�7y%���l����[�G1�b�`�����Ýx23á��+��PzKߖ��J�W�\z�=�W���4��	���Rk�I��;�++�Z'������Vj�	#O}�&�H�,�V����my|��G�2�|�����j�n"s�v:e��u|�θ�7��1%�O=���QP�}���t	��(Y�.*� OW[�����Գ���=�x�IeN� �N�p\懍��A|�%?�������d�@�b6s���4����ʖ#oi����y�6��J��� X�g�z���<��wf,VV���!)��x0��g;�1�-������Ij�c�l�_��!��]����P���*!��5Z&�԰R+�0k��?�)�޺̈́��b��b(���UÔ�8GS��Y!��ٓʥ�]�C�9"5��ͼ���٧��ʪ�ӡ���Y�ɓ�,�2x1�80��|��j��'�[����}z��t�U�7��:#]�{�s���q��������I;i��� ��h�4���HHF���'^��z�A�I�������ώ �7'f�$�'8<�c�
�s��ɟ�ѭ���ߗä����Jev��r���>hz��j��G6i��$�>;�<�n8��%��u�K�hd�[pb����� r0mG�����Cb�����'��4�]A7� |� ����&2 @��	�־�a=�6���LˌQ�"|�vD
�nM[�NI�}���ٖ��v���N���}�7%=##�LnaS�3��������'288t��9xPZ��׼�%��ޓ����C�ӓ7�i��e7I����Ai��Y�󞲰�A��י���8�>=3��-���Z�<~����}�c�q,�b���r���p^8� ��ye����*O�Si��2������13�ADs��ԁ�����1T ӵ�@,w�_Ȧ(��e�	:��㨢e��EOO���f�6g]��7����2��$�-�x��6���xl!�tzq.,,(��,�`����W���C����&x�*6�²t� �7�U�i�#fҮ�1~��"|��l���dAS�֖nk�#�;�������c #�_�cΚ��d�����F�M�ϲf���V��Yw\�5��K�b'�mlt`������ē[����w3��Wx���H�BG�QA#�1�
�ST �.2�b41w���>��g�:JG�"���/��>ϗ��oQ8�4�%āf�K����&�'0ڭNfC�A)_07��:X�g�D�L�.p406a��&��A�E2%v�1����F��-� ��u�D{�-ANn���:��Ɵ�ȌG�9eka[���^%"M�p��JP2�`"���TkQj�,�� ԼOf��Rս�d�h�5� �ͩQ�i()�Sdjl�S��,����e#S�+|9I������_q Nr��Qf��E4�&�}�_?l� �L=�Ji�_ɵ�K}��=<��$���m^����k���?/���`��9��%�?���� Z�1 bM`�+e/)�z���Ҷ��$��^����H� ��P� ����u*�ThLg  8C��|���Iއ��u����Oo���(&��"�)�������}�Q,ȣ���LFЋ��$��^=�.�*+l1[���,��H`� ����7�^�_�P�Ђ��N)S&�g��:+� z�_���t�<�V�����I ��ȁG.\\t����3�����_$\�Q�J!�o ˰�u��Rz�Q o��!ṴX�թ�x@C[X���1$�i��Rd2���D����,���Y ������e.��'ب_��/@�g��O�wr��}�ѹ<����\Ǎ +5=/�ұ�	}�ʫ�_f��eFZ���?B;�����/P�i�ct���w��֫�>V~���?l��3x��Qh���/xhVta���1���b�z���D��y��\A�U���z)qo��ۿs�u�0�-�#T��Ҽɉ�
ɱA�T��G�Þ�1��a ;aˁ�O��y�y����_�j�{�ǠΉ�rsSё���X��|�t�,u�x'�"�=�8��.�O3�]��;^a8㬦���p"�(GI����}�+ա�trQ$�1��;*5 �Ob)}�����A��?�QzN��v�3�:׈m�S�����(�w\�Rb�ڨ0�*�#2�Sn�u ��c(h�������[��Y�l3�Sx�7K>�<;��I�\}��c�3D# �J��0�^� �,cF�8Go��B����.W�ğp�������kҍ���^��K����|/FL����6��q�ߘ&��%�������2>Z~��:�.z��ɿ0�� �;%~*�ka�bW|���Gf�3�0J�\�������#u�p�N���ic��a����L� �"V^rKn�u�dU�Շ^�����փ��泲��.��� 䐰g*Q����;5�F����uB��%C�3��A5:��N��~s؊%]��X4�'8j�{s�	�IsGͥ��V�93DAq6b1  ?bx�c�W�5<�w�<>��;�d{���P=a�3Gd�R���W���`��e5�)��+*^{��n+��(�N���D�f�H$)a���,��!A�Bg�?Qx���_��,o�j���)C}<���=��b*ڔ2'���4X�L�û��{>�a%
퐰�����D!j�9ؑ/�ذaB,�Dh�b�_^����:H�-<�L���v"�t��?��Q��<�~�_N���M���� -"�ȁ� /x��}=t�H^��t�c�Z6u���X�\�R�?�~�ry�	N'c�pC�Q�=}@�89B�v&�/@���k�}C�?c�cױ�AR�vN�m��2���Ԇ	�?s�,�ԓ���+w5@�̩�}�A��T�ߦGŋw�jw��;��d�S��É������1���$��F�0�ɹ�P��b��U%�a�/z���+���  .n���dо��]��l�����m � �9 �g_j��)�)�q^��J=��CL�$`eE�	�q��S`�Pa��!�L��{�:r\5����.��xO2}����z!z���*7l��1�=�����s�%����6�ԇ�� �>(og�c�U� ��>b������\�b
�=.��}?5�J����7}Zڧ�����|:�2���ԾO�,'d�H����و���50FB��l\�b�.a[��u�r�eO���=��P�X^O�M�3؞�"�$�;>����@�wʧr���#�?�t�S���>\��8�����$��tj���Io�3���8�j�JK��G�m��(� ��a�����*�)����m���'��<e�M���{�K�X�i=���:$4G�9�ƴ�X9	k��^,�-�MS�xs�����+q��	P�d�nb%��{2��{�x<�V��5�ۗӵ+�/ hS�E*�ZZ7F�H�;�(x�|����1��!1�9��}�R��ǮKGں֬�A�d�@2���,e
��7��NQB�D�O���*	d��u�a��_ʅ�E��� b� 8�*xFЮ>�3��'�l`���pH!���$R"� ����六�'�8:�OԆ��#޿~}%ɇc�wW�FI�|ɭ(��-~Uo�s���.+@��� �+ɒ�'�1gi������މ�wib��ҏ�L��?�iǓP�������7��6�7n_ƒbV��H��	�N�<�y��+�I���7�b�7�s@�z��׳�Z�!L�� s�<s$ �D����)�<	*+���8�o���@]��V�;2����f�� ;��o�0NU^��'7B�ⴔ�z�mQ��ӗF�h}��1G���>!��^ �j�9e�S��z ��o��d�O�E�[h��K 3U������d�×"x�]���:��i"�ғ�f��WN5�j� [+P�ʊ�Qt��d��� �#7?�I<������rsa�db�`��c�@S�⨄ku��&g��΁��'�-�]JׅWb�W8�$��ơ>���Z�s	���A2��/�����������	��,��dSK�^�5Ϝ�9���30���8$�F��\%�G&���&g�$4�H"]w�������Ɠu�{��E+[I��� ��yB)�c����-�ols`����ö��<1bì�+�])��]x_�+��� ��F����Ť�V�7Ev��:O�&��%��!	��$�)]��E'��)���uK���ɋ�[�ς b�~��U���1�x��8�aD ʒ����w!�%8μ��EqT:��#�P7D�l�T�}����i�8�L�eF{�� =��kn��o�ZI�e2Y�"�:0)�/m+� 3����h�1 ��-Sa���NJ�Φ3݈T�6�R�X� 2�R&}f<��1
��q���}];�8�"��Gq]GM�d���49,��e^���P�*%��TBN�_�(�X�v��ʰ<&4���G��4? <�~����<�JW�x9̒��s�����@�9A�$�k�9H�����f`t �ЗH0n�9+ T�\p*�M�"L;�גG$@�3,Q����Xa]0	��Oa�+z��NlXg��;5zj)���c�~ޱ�=�գ��A��l34��Z�E��=XG�8���w��N�E�Ϭ����m�]/������3�a_BI�+S�(�����<��q���YV��RRI�'�M� F���PI���P@VR��#2螵���Ҭc$�0��F"����Y^Yp9XMC h䚽����c�W/�[�G�݅�`(1�bs�wJ�0��c����(֯�ȬF�-+zP��m��;��e��Τ�a�+���cUF�x���4_4����BC+8��H���~ Z��=HB"m[��
[���(���ڒ������4��e�S-E%z鑩�L�0/�?�\w\߲߄ �&���" ��4	���E��@D�tB�+�P��" MPz�*U��k@頂���}�����|����=;gf��wf�9��{E6��/��6��/�]���s[�����t}_�B�T	T��m�Ȯ<_��/:+Iu�m>��u�W�!2f6��I�7�m������8�.�g�W�>����Ș&ϫo/��)�u��qq�%�L�g�����	C���S��8Fe��b��NG�dƩ@e�8?"���(�>������[�&��)\[�����?��,(K, �$L�v��k�˔�����ŀ��}a���(礑��b3OC����«�vl���{YB��P$Wz��׊��a��
U6��|Ӧ�,Y�D^�~�%U�}���(��|��$����6itY�N�/|��[��=�|?�0>@f��Ѷ�=�;f�w&˛��D
܍��韋kx�%�a0o��� "V�9j�[>m MU�i���W>���2�(��]����܃DJMO��0/����@@X�r3��-t��X&��ia�U�l��<�^@K��,�q�ۭ����Y�0G�/[W�������G���>�k�71� ��B�#<��E��3"r��v��2�Z���z 57�)�I�}e{��[EK|W^�F�(��y�c���B�T�*��~��v(�Tf�Uo|�fz����SǽMI-�^�p��T���|��)��0 X���	o-ڈr8�U��Ƚ���I�����O��TM�%��`!�ԉ�t�n`�6j^�T��J.O�sn�O���{�"˩�L����|�̤�H��/�:��\4�خ������&��OT���&P���˒�6�ٺ(�3�4;�@�t�	7�q?Z�6k�4}���V���M���$��t�*�L��`CS �Q���M�΁)�O{h^a�oa;�g)���q�e/�aL�� o#W��u��S\�0i��5��� ����!�U��u"w���ůwLt�ty��i�T������ɕ��UR,4��'irRU�������#��:��ܒȐ�����W��g<'�������[����Ӥ���F�'� �4�p����~�!���n��|Ţ��N�~[9G�_|0��Ǵ�wh�2!zy4C�AA�`Q�:��(����
Q~�r���l
�o��eu�����/C/���+���*�=I��}��#���o���ݓ#�E�5���
L2����lM��� ��=<Z�	��k���-�ƧbL�p��o8�����g���ߡ�=�p+��9ղ/��%���(����?�O�]�Fl� ��e����l|[�����*W}���!h���Lĸ�(��W�,�%Y�����u�tp41C���B=f I��f����%���۷o+��f�*u��'�����&A�N�Y�Q�)!�����G�u���j�O�J��}��x���
�:����F,]֓�T0���@ Xj-C���t��s̟�*3ͦU�io��Hn��K�q��q��e�x��t�H�y�*R��/3�0h�x �G�[�<���*�@ï=���B�����+Qt#!_���8��ee5��j=��ֹ!�~��L�"�H�1�ԋ�����^���c��ʧa95�E���|�ApL�bKe���	a֤�+���eg�}�K�Rwʋ��d,qXz��c�C�[r���Ka:k,0�_dm�\��
n�[�����,;��CJ��[�k3�]��Hң����~��5��	K�/�^J�=ܪt���^{�ٳݯ�-n��5=d�ĵ�-}y�j0t�ZԮ�*X�]KWӾ�W1����х�uU4���cc}���Q��9�NR]iN|�(С�T�/����Rk�Y��q\�2��=`垠=�2f���D9M�9 ���$XY�p��ہ��RFC9�Fm�۶e�n�ҰZ�K|`D�ѹ8�~&��H�oPR,y��Ch���Ҡ}�;����-_��wo�zp���ng>�i�侒ͱ[u�ulj�߬��a#gӮ��ت@Z.tr� VA!UP���57o�g��g.�*F���c���о9��y��/-ʲ�q��A܅Ӣ�:�Ę�X��Y)S�I�R��������g_W����h)�	v��h��D�;��ɚb�]�w�ӹ�=*k�ߋ��aP2����Dy����$~���a����T���.��Ԗ�'d�~t�����W��>��3f'}OS����<�� !U]3]���zhKT�J��04�v�o��3����-�?ʽ��$��2�,aؿ|�X�2�Z��^l_p��[D��&
4=[�������d�[���?�7J(&qt3��+����o��XMу!����?�tHxoY��ȃi�W0�r��'ұH����м
�M�z�=���2L>	[�4��}s,+|\�I[]�[�*��h�:��`0X��G��".U9[��b����̦-����
��oJ�4}r�Q*�ݙ`U�����ќ
�oj7�|���9���ZY����@��qƭ͎;@�$�j@r���+�?~�6�
2[x��X
�s�}۠sk�=�"�	���*&>�U��kzuѾ�6p���Yl��x����,����>�g�E�
�M�N�Z�{�������}x<�xrMԬ*���LY�ҫ��������0^y���N�J�ޣU�bR�>�
�b�����t�t��72���DV��g K��Ed 6����uA���;���R��t��_�Q�3?�N��ԥ��M9�C���k�Ʌ��@������¼��Հ���tWP�P)����/LhkkS@4��-A��w6wd}�w$.#� ��
-�L=������0+[0׵��{��͹�<�dl,~����������s0�|��n�rX�'1҅?<��nsm��)�R^��z����=\��j�F8O�t��d�;1�=(����F;�h2���@GK��5������Y�{���ѫ���G�*�_�$;C��Ս�N"�YO��
0l�@�ض?�P��3k�{����	v4U��f੼9�`	X�"����Rߺw?	�ڝE_�*�>�X^��7������'���B�X��*�<$)��O�-������]H�Z]�[Z|�
���ft��� �� �<��qd!�����*��6CQ�o2+��a�5vt��p� ex�o/��}.�)�LT�X;w��5�����]�y�o����K�r�A %d��@�/��L!L#�u�Vs���eE��L$���I���w�c�W�*���f��c��@�9s�\8�M�9�k_EPɇ���:ۥ�_.��hI�Ϋƶ,ә[."t<��R�'e���q�jɴ%��aؾ�H&<yᕢ���s��[��iWdB^�L�~##���]c��8��i��Φ�;���K��ev���Y݄�o3Yd�J����@z��ͳ~l@�p){��,,-ͫ��YT\L	4��4�_cǤ$��ks9���&�IW.��W�ĠwdY@���Jɳ��7�����j�`xR&z��O<?kB�}��\ȶ#&qwt����y�M�QH<h�ؾE�}+�e|�*�iPzb��:�2�g�C������_� �8�;���U�����2���k���.�+}vt3���S��)��{�ZY|yp��wI=���S`��J���XTQ�xm���X:j�������0����_^�)4�|�`g)���9�-�tgz�]�,���Tm�Q���e���5�_�[�{mLjh:�G��,�E�Z���b�]!���4Bq�����K��H4al��p
4�G��8���H�������u�U�)��D˰�Z�!���Xdݺݸ�"�$=��#��u�W�F/����F�r�D[��M��0�;��4�Yd��Y+��*AZX��n����3�S��������$�����r�prO���& G=��k.��l�V��|�5�Ԯ��w�ߟC��1����0��]��7���'W���g�uk�*������
4f��Z���/�����`H;�u)�B��47�$D����ܱh�G=С 1�z�W�;r�����Ȇ=Z=1��^���C�lK���S�f3Ǘ�_ɢ����05�i�H�U��F�|_����$��}ƌ(���k�0��|��z��q�+ߍ�V��­�Pq�����~|g�ڡ ��G�8į�l�f_����Q��Iɓ�)�S��׀~"Z�<�ڏS���ɓ+U��4ws���njo���,��c�&�{�W��1xH!�Ʊ&�����TB����MO��Ό�z��\��e�t<,�P #��x�l;��7jcq'���y����3�ym[C(�~y�)����!�x�S$�?�l�\dlB���Y�o���NEw�?�j�п�1��U�$�G������e�y� ��.y�u��Z��'�mk(���s������Ʊ�(.��75�T����i���%c�Ю����*�d�TޟX�̜�G6�����L�7;����A������8j�Wr"W�O���$�1�<OU�:eTQ��|^�f?�����6�[�
<$�;FFC�D���e�uO���+���־ko;�>E���H��m��!eh���c�c������5���� \��sc�����H��B*{Xy0�MA�N:��k�����*������6����1�Z�S�f}8��j���i塸:0p���*�}���'���E`�+�?�6 x'-�*`%�TP� pr�FHpA�C�X�tiX/h�go�W��Qy�@d�����OM$3���v�d$h� ��}�3:�M��=D
��9 ������/�?���R(���#���ЂMԲ�Q@V��	B�d(���<��O�L�ξ�P~����3x�Y8x�� T��c?��r�=,(|������Y,5'x>��@�졈�o��x��	��ʌ��: H~zh#�
W�"������%�=S��
ݙ|��,���\9{܊��Jfx���6$��E���݀���yk8�?Ӑ�p��C���L�z�p�gC	J��S��ɯ��9]d^�1� Y�{�<k�>�����!h������\��!zl*�WO�ϓ�SXl��	�ߊϡZjz�o����PK   �a7YN�v4	� m� /   images/4949577a-1080-4c93-a0f7-9bc81c12f32a.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   �c7Yd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �c7Y�]��N � /   images/907530ff-a8af-4c9a-ad67-f4101e76dea0.png\�<���?�m7vk���Flڭf�e�!�]�m5���J%���ӧ�P�l��˖��\"�k%��E����0Hc�����������*3����y��9�׸q����/v~!$$��_�)BB�K�����l��t�5}�>��;-_A"�E��?��Ղ*$$������iS��7�g�M��{��y9	�h4ŋn.T�sN��^��xZ;���:���i�������`�RaGo������oޭ=&�����O��)�ʓc#ʓo4B���&�*��.���C�7l�|�돯��b�z����+��^��kY����зR�k�f��IB��>&"↼y�G1Y-nG�W�m����)����}CVܔ�������I�
;nX��r����K��}��	VYN#����� ���V/��)k���rG��]c6���h��S�T}�CV�)Ly����Z�li�Y_��ū��n^���LL�JH��t�3�h�=+gfR�g�n��k�^^*�0�K�����W2R.hɘ�,3�8�K_ZY�&_,cqO��mW�!'(2�:,I�1:嵆�����^��S��I�������[���^�]�Sq��K&��$M'�IVi-��ۧ��)Z�w��C���w��7����o���>��~�z<���h[[�aZ�z�7��0��.�6������AW�x�z+#U�v��\��ڵ�iܲlzk��Vobbb�J��������$jp��0v����K\Y�+7n��S�1�4{;��1�r̒{�Ai���o��z��U&��Kq�,�<O9�򱪴���Ɡ�x��_7A�������TU��s�k<Ե����)��Gs�)�p�l��U����_{1�58�
;�譓���y�>ۈ�j|�MjBB���i<j���Qe>,�6�h����dУ�mh��E�Q�����Uޕm�S�#Jb�U�����ըL���賫��2����O�h�M<b���%MtW>�njjڣ��#��	���.�A?/�P�o�(��(׻�����Ǡ����?��*����Kݣ4�4í��)����I߈��6�^#�߾}k��QW��X��4����H��9�FwN��~m�%7*i���4��e��5i�X���]_����G7v�L�����JP9T�1�s%���b��A:�k�\�HR�]J�~���X�,�<`n�]vG0��+놴�x~}��D7x8[<����=ޔ�D6�0�#�f�?;$����*]LMMYѻ4!�d����E�_�e��-lmul�	'H�
�7��F��}d�+4B��U>=���]�>�o]48�\kK�kva���zյt�7�&�0�!���ۢfôs�^����)]|zk������I�*�<L$K6��|w�מ���<��F�ݍ��()5��ώ̽�x����g�2�27���a&w��LG��a��N��p�ܪ:�Ru�)��Hw;\��I��%_��8���8�hڳb�A�>R���4w-**jϋ���S)��\�O����)T�3D=��#����d���t8�Ӝ*[�g�SZ_��������b����7��z�Z�o˾�/�gxv<��ܵ�^"99�����Ѻԃ�0!F��&�k�����m�K��{�L��߸��V�).ٹq�S�TaG�m.��͍��=���R!6�{-��%�f�Ҋp�tAs�%x�oZ�N�-��N2����ݻ`W�"~�������N��E%WV��N�$�D����ip\H��0-�����,u��/[f}�ڂ�[J�2�!A9e'�	&$mi�zK����p��Ǳ�3���B� ���r���F=%��ꐠ�����\=�������9x�o[ )���tE��Ǐ�,M���МL{�JǏo����Pg��f�'`��6�٤��mMH6ゥ89�Ǳ6)΅]����������{���x�<6@ou�s�����԰{��V������~�*ی+ X!��ge�?t�޽����.�i�� �{1_P���ޞ��s����.�?�z3"���7��,��# �6�GBh�1�,!��<�UU��7�����W'�+�5�4�q�$1�ꗖ�4c#���&K��s��<�
O����e�l�����G�·�?+��t)�a��FżO��31�2�w)�Gk[�?~~}J��)��\\\Ģ���1�I��!������)�忸e���1%M�ͫ��Y�M����������1�h�,���&h�����n!ebBweI����cF�dc�]��^k�x1���+I�F@ȓ]ߠ�,�*
����t��2^K�lPv����{R��a�K�� �T�R��&d�O�{噽��K�g����v�Byv�I��/)/���V�٥�nX
����������cY�`h�r�n-�\�WG�A�.:����� |]B�
�g�N��?�T;tHf��gM{b�}�hzir�����]>=b;v�8d%��r;O<�e��#�z�l��!q�v���N�S�Hq:��rp����<�����f:%�}���F��0myN��\H<%`䮹����,�~}ST��g�uu���Ϻ����,'s\����"_$1>����h��>ڻ��Ł�����I�"�Z��}>=򳳳qTf�al�O��K����
�qp��'�Ѳs��$TaZLe�Ҩ��)��Is+�يx:�Ǘ�{�Ոx�-�bk��{*2����&��4�dHb0���r��=�`(���D��ӧ���W��kݦ,���}"4WEi�%>Sy��u�e=���u��}i޻o_��2^fҬca�-w��}_�~F��<�g������gΜ������C�^�6)5�:	�K,I�H\?��������vN	B��e/�'�u~��dQ�}j�j�J����*���ڼ_.k��꾵��+m�-L������<v�`Ne�9;J)N���F/g�oP�ٰ�ߖ	��t�Ѩ�)�t@A�2�P)�0����ô�u[�A���K�?�m*�#�@�M�Ux��ͼU��;q����1�\[��B�@��Y��o\��H�؎���0��#Ii�K�g"G'�{��U=�h�Cv���PM7x�6u5.���ܹ
��,�� �\������4sብK.Y�Xx���%J����ĕĩy3����S�o�{1�c�u|�q/�<l���8���1Ӝ��c�#^=z��'�R��1i�e��<�]�%�9�"!t����Mp|g�6syL�e�\g�s���2iv3�JU�$�(��^7�:�����t:u�l6�Nh�z�<�$>��'�ϑ�*���u��ŋ�.�!1bj:�����r��;$$r�x�O��3�؏��c��|�)�������L1+��%�}���\�����1>�D��t����US�s�7�y�����*K}O�[�Y>* Aa6��4蚘������G�9So�`	�3�ʸUL���a��bN��ρcI��C�_ZO]]�m�c��m�mف`y/����s���q�#���y�����H#{H�}.ٕ�_�.� �����h�D �l1]�8''�F����n2r���Lz�A�������2��#��L�M�����;&!h�����$��$%##��o޼�B���%�_�h�c����2��O��>C/O��"[�I�� �@W���w��k��RJ�>S��K6���b����H��!6�=�>���������<��N�7D���LI���L�Q��?��",VRNXl>3��˅�esC���^k��p�MlX��h�D����
�Dl8Iג�𛾴{�d
*KM�*5؝XAA�UbU�u�R'�x�pa=�	*�zu:d$ɜB�KIM]sc�#��i����7"2����F�R���)z�y`;��K�w�
O\�<����Nu��""l�>�+qO�����Iԧn����0�|!'����
*�T�C-<���a��yDbLA(��j�c�J� 2�ܟ��ݟdbB�0��|����48���w�;l]�e��%/��������#�����?�q�R��g�-C��H�m��V= �������PmO����=Ω�����	}�ɐ{�&�%�qa����赹�P�!�R���˼G�{N
;/��<��Ď��am�a��]J�2�(��e��aB��^y�]ys�������h�KPQoG�X�K���]���1a/~��b5�� ��Z>����'� 0|q�S��ۉm(y�FM���8�������pI�mh�ak8_���$%-��f�\^�����o�UJ+*��H#�=�W�Nj���cr��$F���BE��$���܀�5���;��4H���'NOB	`NȂ���ƿ\�������XȌ��+��e�v�֧Gě�kC�L�z����`0J333���dr�m$I$�����ǚ�މ��p���W���� �ڊ�����g�ӓ�����R1��� c"���k}I#�uC3Ő��b@uf�ͻ�>;77���E��x�s��Z���Pc&k
�{H&�Я�nddęL��C�M�7.}�I��K�DTh^�,Uc��<��LK.U\�������,p��]�['o_z
oW�,[�5���~Jd��x���Q�m��<WK������&	�O�BY���ӳ����"¦W�䭴!���G&I�ۻ�����#��}����	�_;���bZ��bI�ʒ[DG�t{|z��qx���� f93�J[�P-�oK�i�{��俠ĹQ��w�`yaA�d_� �N)SVS+~K�඾�;hyR�*�U�M��d�#L��'��?� ��ԁdw7DU.��f2h60�nY�u��ݎ�jS��CU,�?2ݵXW]7N��~�5Ч]br�n~%a�{������PW��c'��KߒIJP�B�e�]8��XM����3�溱��lK�m�_�
Wۆ���M�� +B<�<a!~[��\02˧' �l�V/��nݺE#XgY󔽉��U�Sn��~m�nX2j�1>f�Bm���)"i]bv���%��֪:%ޟC�Ҕ[�[�[[�#JP���sRo�AE���{�B����G�/�fՉX�%V��fQi�B�U���0B1хqH��Q����b0����ej���- 12�I���jH�x���bJ`��nc���{~@�1��T�h�@��J�Zh�)jY�s(�Y͓��w���;jp��-�
Qtv�G[D[`%�7y�k�vuu�v�e2��ϑHM��d���qq����	LH5������.�q��"�~#n�@����'��}v������;d���P�X(.n�P)�}�E��TВ+�o�QUU^YS\���Gh��UN<x��x�[�������!��t�b��~�[I�����8`S�BLu�Dk�����BC��j�na�}�7�T��f����0$�Q�'���ږm�����!}�|HȪ&8��&���	.|���7u��3��1K���ŚJ�̯5B/��x��B��(�98�������1��R)P��c킔��ebl������Kv���B=쪟tu��@_pd58[�j[[ۚa6 ��d�Sb�é���
~��f�8%;����g|���ʙ����ՑU��	|E��snDTTU�ޞ�[���ñ�����RSSS��Sgb�����6�����4°���4$�pWG�	�./����T(���S��م:qI?!��'	���gϖy�C�����!9�V�I%�rg�!Y��:��^������`0�+���%w*�~�
�(Om$)\��^���q��@Pb	[z�]�Wo�o�u��Ԟ�4�NY��\}MESs��N/�C��
�V�eH��ܒYi'�(R<�l����N���I�;��}�a���;`�pb1��x1��qw�J�;Z��-48\�s1��~��?'6ӹ�Z查U1�U�'$��F�0L�����i���"�Ɗm�s�1���پ�n�p�C�/0��la�YR��I��^^�MR�J�xd�)�h�:Š��$�N�n�{��Io�RS���K'	�HYz��b���Vm��z�8�t|�d���\M�ޏ�׌�>�mM��s"� �ݤYy�|���*5od���]����I��v�Cm�1w	������imm�_�V^�cf=��W���g�b�Cs�K�)ZH���������Kh�}H�*�˛f��-������_�s����B��d� �<F9O	E'o���5Մj	4�	t�g��C�,�Ǉ������{�s��GbccG��ӫ$�g����^i�Pȡ��QP� r[ab8ͅ��v��%�.��	�	�8�A��$�� .�0;�	C���Y�[�_(uX�""�pN]m�'r�nc�MP�uזk�N��u9��j�y+�%;�,b�q��N�,�`��z����2a���$�=JEX��Wyt�Be��P3�e�&��÷۱��dKD��m��F(k������4�1�L�W4bQJ8d�v)ʥC��\�n�~jdj�P,��j�J"�^XeC-�H2�J�_��]���)Y���)U~l5oN��%x/0�X���@�Ν;v�Z�.�Udv�xJ�bmmmj����R'�W|��nag��&��-j���+�%s 2k��);�
v��?w�������~F����!�8jU"u� ��������{u{��gQ�G��L�MY\��Yh��Y(=�����z���g���G���7��$����%��y@�T��h�u��^�r8*�p�+G���*55A�?�)'-�Y�8�=�R�a�2IMZ���>��k����^��ӓ糭&���W�9��kam]х��$��ĠV�h���\�FaQ�����ur�X��1�CR��������I*6%�Y�=;�K �K��~������Eз49B��V����Ntr�x}�ZY>��/
s�eK�"yv#Iv����D�#:�ؙ# ��2�;�	�޼	�����X����b(Ƭ�\X���x�լ�hr�9�7oV*EH&<����ޞq)�:��>C��-i�FFF
���
��#��\��Q�����v��	�G­�j%��oxe0�0MMM���e/�+5�^�������v�e21���C� �,����nk��������]o݇N...1>6��~"H/5�[�cBFmג,�y�Z2}��x�sss�fD��H#S���T���������)��7�e��gI�^�F���)		��T��ߋ�X�C3hî�ҶQ-+��:_v@M�������atnoI}��J{�[9���2��(��룃���R/��*����[�(��#�����9ZƤ`lR�(�l"�,mw�X ��!��ۯ$Ƌp1]m�}nt�6V���([���$\q�]����ƈJ�O��3N�#��S��r�E,t�E����r�%���~gt����#�:�ʆ����+�eQ����
;�a��H�Z,�%;�j,�k� �����:H0�rEu��ƶ�d���+7��f�/�|������<�����b*�in^��*N�J�'QK��?��6]UzkI[lS� ��9�|H����h�9-�;Y�p��Z2�E��\�-�oj�Ֆa�[���DH�^\S�T9������߾}�"[�k���
q=�������~m	D��T�v�j��7	�.d�%P�@&;Y��9�dQ��4���I1�D�Rv!�ц�
���e��U[���Z��AQ{�-����!9�Kʒ˿d�`���,	��Ҝ+��%8���<�V���͒sx[�y?���_I+Ÿ����-n���l=@�sPSx��VBBBs%݊�v��� @��/��3l�4�FGG�b�s�(oǠ�����;.���$*���Oe�K�ٚ�Y����E��:;B��I����Ҋ�����&�P��B*?�9���\�ijrJJH�O�h+T������䖝�~VnO��CY��=50��!J��]������>ZZ�T���_�1�(�եEa�Ɏ_���H߃�X�Ш���0;���t^Z�Կ]�݌����N`�H
�tJ�O�1��-�΍ַ����TX���:3��+	yj�8��T֙3g��髦�o�Qd��R�F�gI��[�1�e���k��*~nRtb'��l�<��P�-6mK,����[�����+�4�dn�m�La�a-�SǫɹM9!X�I"���l.��R�����R����X����KLL��~E�֜�pӒ�>$-j>�.-�)n��(Qg��
ǹwj�����i0ߚ�~�i!�������T��q>Ѕ@hI.)��������� W�5��mC��!�M���19�M��N=�����ļ��WYYyXZT-��ʮ�n ���\�	J�i�a�8��l�Tm�r���$�����������#��-�֪�¾�f�l^mħ;X{��1�E��.{e��.+i~��*�zA��"�;ˍ�pPZTBe����ˠ?���3ɩ ����Ą�%\�֤�y0tY�1��cWV��'��<Im�4����:i@�C�f���A���a΄{"R����b��,����ו�ħ`mF��o������Es�X��Xfd�q~��+>%D���f�@��*�T8�.����4>�/ضm8~�U�S�!�]Ju.E1'c��Z�Z\|�����!��F&�
���TD<8~z���������)�m �����D��o���_�����me��|��ݞ�[$'�c��ܤ�&����`��1�]��ɈW\�Vx#�7���<Ls1���$K<{��s�ja֓��rqq���X�\�5�Kb�.�^��#/�/��K�8F�^s�>�i��O�4֩�ޚ\����i��*v]�ܝ��HR�Q��k]^^��<L��}���qP=�V�~�E�d�+�%�P�=�0֔�)d���b���t<���- [dEv_c`WH����(�t� �\X}��_�E�q�N��4���w�SL����33~�J][)��NE���lX����֧���ws����șM=�m�,�Z~6>>�0籌B�n�%K�9(aJ��+: �uO���}�.v��c����gϞ�D��܇y�s��RYի�&:��)Gͦ!�W����ڡC�)�ű�T��T�mT*՝��,��h�700��Q]�eFa��|V`e/�ZcQO���,5�rN�O����ڞ�D$��WVj���V�i{�$��*���V���2j�I��[�g�-zh$aj�q����q<�'��a���
�Q��e%6�<���Ȗ���ac�vP�40,�Bc����gmlV(<
чp6�����!/}�$93�<�����\�df)+X��m�d��z����n{�m0|.a��
����	�m�g�v�|�tg�u� �@���T�-�@V*u4w��΃M�41垬� �kӚ��]M�5-�҈5��$E���[NU{Ѷ�����!!�w����A��]���W�r��Bm�'�3f_/MU�y��Al�����z�sÛ��mE'n�{RR2_�Uom��KIZ��wh�k�!XNpC�e
ym�M�jh"v���EEs7�rt�;&�u����q�t�˯�h��⯬��:�61�!�u�0�ecQ�RDć
B�	i�����xGNW�����'�פ� �hZK�aZ��H�ކ�ZV�b���H%{7���O�qR����n*%�ڧ�(��k(S��<��:�1����b�9���a����D�P��7m��^�c[����[.|����������;�tO��}R���W��}4ͥ�1�y��6�e1�攕Y�v!#�vF>T�� �Э��Èև�{z�L��(����X�a��U[o7h��hT��9'6.n�j�B�����q�?8;F��}E�r8vm��v)�WǶ9J�������1"���kn�w�{N ���;����U�}�����*)����&�<��� ������mܵ���\<7�N�q��.\T�8C0�疭�H]��a���[XZ��D��ș��.,���3��U�!y�b,�� ,Z��@�;"RM��r���t��XFV�8���F��QJ��CK�ߤ���W�6�
]��&Da�	��)��
�Rh���`�u=wn��dc�e�ht���-�Pgw�)��*=�T��z���>�&�
�|��H�����A�O��]WBւ��Bh��21��}}k�m_�Uj~���!��ݻ}���į���.TS���d�|�/��n�)�T_t�̼��e��Z�&���� ��{e��>��W8��y�?:pq,C�֭[�
7۱yd����ҽ�|����n�i��P}T��0��ȹ�����<vi#aii�ҧ�tO���Z�@��������6�/�����I�
r�����|�{E�k+�TN���pyW��:3�rĭx���zy��	T�? ����L{��܅��s���#�Sx2���w?|�����!����bA�\.7f���3z��ҨOy���/�|�Cd XH	�rd�߻��o}n�Dh�B#f;���<�m�>v�+���1?�,�MO��ϘB����C�Â����B��@�쬬�r�GqAZ[P���5��^WW�w�T��g�����iYY/ٻ��^JB���n.r�rV?ڐ_q&v�=��ck��+q���8��!�ؑ��� e4�G �Hvҷ\V#��Ei�<�;^sS����0���E�*�9���"t�6�kwC�7�Pa*a��ɾ ��J�Ϳ �5sP���K�&����Z��_��T��x<]�Ffw���SPV�h�d��y�L��iTT�!]'��EE!D� �=|M�^�F�3�3Z2v�����E�.���k9�xc�E�6���@㇕��ǀ��رcGo�7s�f�7?"�t�^��2���Y��A����%��qZ�*oS�#��o=�İ�!�6�����5��÷>� |�CIpD��34���#�㦩Yv+��k�-�P6+)ˑ@Y�.�"t��k�YY!ܷ����yg1��_Q�����do���c��k@�r�����#��*�g�x����(��!��X ��I@v1T1��?�v�|Q�`
�,#�7��s�ң�Nw��`~��鉶�����&�V�D�Ξ��q$1���tQ��bs�2̞�#��8�Q�M����}s��7C?~�,�ɇ�v���{�$"e�I|l(A/�+H�5�0���H%*�����i�"Tpk�YпԓR�������y�*�qm�wC����V�/�~Wߔ�^�Dχl������+k��h�H3њ�=�Ն���;�m;�8��"vJIk�'B5O��>��r�F�����roo/+1��>vUVV�C��y(t1Ȕ�ТTb)?�X�>��/�1R���M����C�A��~�IU��N)U?��IU��0E��w�0-~�I;�G��Ht�����D	�ZM�X'UՂ|�@)ׯ_��\4���[c#���w��8zp�(�=�@���߭:��6bO���� ~L N�$x��o��u5��Xq��"�f�i�q�<ޕ>
���y)a�.��K��"(����܏+��uKE��nbj*�K�P�⵿�^Yٽ��j��R?
BaJ�根)y��n�m�		��;ru~��ч� q�d;�7�+p^sƞ
�����ɟhҪS�<��3Pc]�]��"H���,�����y�]l�0I]Mc�&�������2�6�5U%$$lC-Cg�h�>h�M]�r���]��"��W2��*�'��{����k��S�f��>������#����q����%��&P������v��j�q�m8���t��A6�1	�ȣ$0�k� � uL�QKR4�OZ4<�����O���)An)��Wq!�璣�P�J]��%�v�g��~f��@'�Ҏm֚���]�Z��%$�3:}roȗAm���oP�L�H~S��*��ATUBowHMM�=A!��
�sI��&6=tש�v��}g����՘�w�^�g
Y7���ɢ*����Sw�c_JA!����!RJ��5��prhp_�����Ss�;T�ަ|a�c��P�ڇ���8Ek!g�s=���n�X��\Yi�� aC��+��K��3vX�x�����@b %�C㇟p(�9��v�5�0��i	Is�c�5(ot<��f6a֪ǧ5t,{PalL�&�c	RTHu��k%M�6�&&�To�,��W��v�[*&�hy�)��C������)���>6		��h���C�)��� �AB?g�J��[�#G�����Կ�&s�$M�Ѣs@�U�]���g�ቶ�J<^H!	�ͻ��Z�!/g`_I�����[`��y�&7�n<��)z��e=���5szgL}3$���-��׷�X����	�u@�'n);LL
]�\Nm��4�y�N�D�"Ӏq���5x\tZ��V��@u�N�"���o�w�����]4�K�_�C�n�~�$��C��G��w�{0M聺��N�V�>�
FH]�����G��U��@L�A�22��*�e��a߼y��ٳ~O�X�S�^#�TTI;�k�!��@�¬,�7�q�Q����.AR���Q�75��--�2}h�3�Ɏj��prC����N��	;���^j5������j=8�Ϛ�+���`�PȊ�?EG2x{;�9J��+9i;(���7D?*�1QRP�Ґ�"�C�5�k�C�r�K����u�OB�)�N�������3I��Ê�X�W�oA��j��*5�a�����D&9��g@M�����V�1>��¿�zHu�,/��/y�u	e�I0fL����M5�˗�����=��_�e([YY�^Nݳޠ
e`
���Ƽ@�f�����W�˚�N�A!��j#P[ͧ��������`	�8@�8���|f?=O�ޕ!������&1=Oe�?�YsI��%����C3�_򔯌��T�,
�k/b����Rg�v��r�Ip�;x��*�pr;��\����I�M ��GyB!y�s&y�U����V�%?U�I��;��3�E<	�nnUL<�&�:�R�0ٜ.28p�E\�/;Hs70�pfF
�G���/���=��ZM����J�M���};%���\�s�v���\y�������;(c���7�w���*$��>�����֢�[0�=S���8�����2�TtJJK���=�i�W��W���F����!)����%��峸�O��L��MLZM�N��(�_7|O�F�n.6+�W���4�L&�I���N��͢X����"�,ɪy�{J�E��Qlc�R����d1ؾ-� !�c�@mZBI�\�m�f���7�G��Nه�Y5��@�!L�{r�K%��ǮVi���- j�	���%�Q�
A��D��ֈ�
;��%1T�tM*m78���(��߻ F�3~At͍%_:Y�4�������^pi`I�JU��Ϻ$��_(i<t��6�哑-���a>h�zI�M�87+k|ѽ���'�<�/�+I��'3�M�p8�I�ڑ/P# }�����)�(��(D;jkP��pc۾ޟTU�7�UZ^�%��0��}�3|=\��`��i�9�Zt|��-쁈̬K��7h[ ���
jN��&��)٭�$�~�F0�'���5��}ȐI�f/P�V���q��D�� �<g����)�,_������w�
�9H����E�?!4DgI�Ez&�4��,��l��ٲIBo��/=_A���s�:�wcT�)f����o�E����Z�:���;h���D�����KlYN 8b�qR����WHc�����J��98Db#�V�}q�F����w�%�K���<j+=K� �<�k��f����(���h�{�#�VU]	Y�Bұ"++���q��d_~U�ڵt α�c�SmЧ��| ��e���9��P��Z��W�2=���*��DaE;���$�����h���H����j%��~6&|y�]�܁ۚF�[�$�lCW����*��&�-�\���K�,W�	Έ�ה�� �ݲ�?�&����ҴKQ����G�+��{���#��XuL�N�z֖V��xIk�p8���;�G�� �B��5��N-��J�6>6Jü+i���S�yh#h����l!
+>��(Ƞ�z���(l�bfFss����_�w�ٙC�`!p�&X
��ZsS�����աV�F�)���茏��)�K�8i���[b�T1�\��vY%�tS�MW7�Z3Y���t�:�φ��Aho����UMi��k�؀�~��������
֭��]G�R�A�p��V�N�S�?�����e��\ mŻ�}u%��]�͐��KAy
촘���X�������R)�h�����Wz �z�6�G$B��ԐFe?�S���</�UrR�$�C��kL�o�%N]ۺ	A�q�?��?/tuy��vH������t8����=�k%����]]ށ����xf�yt�d������'}M���P��'�:kɬ�@iʚ:-!T��)�`)d�Ql�k�H�̋�+��N�g������	V���3�	%l�=���99�W�>73��#���:;�|�9���|a�P�T��)��)HD��:��0GƹMI$A���5*�v�8�<RWW'lJv��i�íz-\>S���#����^~}���2����?�9���Y9�����O]�8{�s��=���Ͼ���F_��"���-��P��ySS�M����b�w�=�(ľ��� MX����Ɗ��1�a4���G�L��*�q<Nqś<�`x���~�ώܺuk*��XU�\P6;;�{
�**Ts��`���=׷�O�w����ѷ?��&�/�.C�[5�����ZY���z����B��J۩ۃ2�ON�*���Uz������Ûw_������!?�u��6�:���7c��"�s?���+onk��{܁���ʏ� ?^S.a�V�p��8ӕ��`�?�*G#���I�Ckk��x�-am��QT{� ���;a���+�'ږ+%�D���q�c���G��Ro�/MOLL\*�wOݦ\2%w�����@�V��B$��X�J�S�������N{����/�|0�x^�մvC�c�;dVxٓ�m��T�oKB5�yb��
m���PWE�?���������U�G���R��G��08���<��Y� 1�SPP�dZ���V��l����z"�&(�P��:x���prr������Mrn�������(=&@&��:*kB�'�ee@��l���e^��w���ڲ)&�i,RX��i��d`f��Y0H=�oG�y��Գvv��< ��}0�c��`��#�SF�~_�J�L9�^8VV�"��@�柠6ɉ�-�E=�1�
��O ����R�7��Z�=���H�������>�bWW�΃'f�$����'�̴�j��uh��]}}k]��GT]o%r?>!A�ݤos�O��k'G�>I7�.R�����<����d�v�i��.��cj6��$�gɤ&e�/���o�x905�F���.//���:j��8S��[{���R��@R����b���U�;]Gܮ\ܮw�H���ǋ�H�޼��t#]�7�Y��.BG�Ð�Н�񄄄�N|���\�n��&c������m.�
^�07k����<��|���-��[*�#׆|i`��
����q������4�9���n������埽��T�
�r�5eؒ�^_��P�kw4b��o!��ÖtA����J?�v����Qv������+q�LR*n#�wc���R?�@�T`�Wg�������	oF�PN��l�?R�p��xY՚H�=Q����၁�&�	n��}׵�E�FMTs.t�=��C���ev�B�����.�00��;���' ��KNN΅�I���f~@�*l�Z�:�-u��T�q
=@�lto���:5���;&�0m�l'@�	�md``��� �����������SS����k��j��N�Nnb	�ae��E��a�L&��E��g��1>~LPu)V8�(���i`�9��e~~�1r2��2���R�2ۆ/���m���������Y 6�q�2���������h�()(�}Y�j�J�;-�C������p��~�e�*풖^�#9�-m��κ�|[	������:j�{zV�f�*�K?c�*�P�
��D���N���x��N�f�هYY�ֶ��wp�S7s�oٹ�S����7�`�[3�d��"���˥ۗ���6v3�a]�ͥ尸�J7��_T!p���Wx�S���/���߃��A� ߴ�~�~���Ļ�ꎢ�R��J֤/n.n�S�5>��x������)���%6N�T�5��׷>������[���v�Z����~:43_,���7���\�gc{���\���l�zc޼yc��x�L�`ȅFH!b��A&�z��-���:<I��O( i�f�&�ʮ�+�������8�7^@E�3j]:F��,)�\�w/++����L
��g�RySSv��Gp{)��>�M�n���ra����g�Th��z�����p�2��'vs��Q���( ��]
�4��@�K`T&��,=�/,�q�̬=!9Y�o�[f��^!�Z�!��D�P��"�9�e@0ʨ#��8;[�����q�.Ģ�x���r��ZIC�w(�`T\Tp L@�_�e�;������,��RS�A=%x4��6�� ��UGG��7z��Ϋ!7����(r�^��Η���従$j���@5a�s���89��%�VE���u]vϵ�v���o���������m*|�|��@
%�\��ɹ�s����֖�I��#���ۏ�
E�2�( Mo�;����{�֢ٓI��ɹ��	ߴ�]HLc��kT#H��_��X,j����pQ=�h�:^j}s�c>�����%q�e<P��!�Nm7C�*���7�M��ǎ���-�F���Hz����O�|X��i����?�]X��%Ĉ/!�B�{��D��f�Ft�G]Zt-����o��)4�(()A�|��Ԝ&���*U`r�]'����Ꜷ�y�F��/����(L�gtT���\��o�yxU3~A�Bc�����	����^��Ǘ���=��*�i���7o�PB�k��zY������5%�O���UmcZ��ޏ�9���8cTe�+�~m0#��ѣ%X��N�a+++wu��K�����)A�\@e���nZ�g���B)5��f��[6�9f+4*�$E,������V�����6�h�]��\2��G
�e7� ��}���\ݓ�_����=�b�*A�u�\�Ţ�����k��İc'c�����d�y�^���#=K�˗�����de�z��/�qP--�ǿd�k���?����f�Y ;�o]�n� ^C�S�.�3�����s����z��]�N��qMt`��� 1x����7TRz>a���ru_�⎛O!�\o�����B����h΃D/w�o��l����`*x78�>�"6���f�(���/�.�^[rfHӳ�3#	��
�X�B�hgX>��*SXz�|x	d�q��ͭzj41���B��zIS �A'�"ץ�M�%&�T���1�d��(v(�#���>�*��E+�r[�REH�q*wʅK��bb�n��*����c��:ǼW{�{z���jf컗�o��grK�8�# �ͺl퀡���_�I|"���̬	U�Ƭ��H�r톲r"(]��[qC\�&���_ x�s��t���h�Bd��P��8'�Nz�P�=��|U�B��om��U����^xx|W+:1U6��-�S>ഏ��>�A���N0�mT�K_���f�[mM�~ff�J�J~������*҄�j��P���ļ�����I"j=�HK[7��d���C}-��_��!ȮBR� ���1�� X��^���� `a �o��P�����FC�a�vY�T# �h�Glնa�'w����^"�Qӂ�tё08��×M�3G!aGBJ�Ȏ��ǔTz����GxrK<�Njj�������ȹ��?�V�ppq��㩂�Dw�+�>���'O�m�Y"���҅��C.�8��ff�P��PUUUj�y�,�Ȯ��s�*rE�d���7��������R��Ӳ����e��^�S㜛S�M���������5ϟ��L:�4o�1��&ж�(�鍉�8	���� ���ҽ�!?`�~�ay||ܝ�Z����r�G�e���vF����w�������_��p��Ѫ�,�}���v��[���ŋ���}�Q�
7D�?X�cf�X��K��J	m?
	}[���n=��u_�+��;���6�@Iǅ������-��x������@� ��9�Bd�r:��]�t\���u�e3�5���������7�ͺ�,~0 U$���TH� �{.�����;t�R�Yx��Eitr�����ߡ|������5�l��CzCV���h�;r�w_d�T\��Dڶ��ۨ@��Iuu�X]�Ԛ+�S�Uh�<��G�>�g�V��!҉<6��n|��h�Ľ��
Zp��n����}\ZQ�w*�P7�����\+���$a��,�s6�Kyk�q��
@�������_V������ˌ$�R ��)���kHj�$�+���q�d���پMW�9"���	ʟ���ǵ���E���J� q�+�~�X*�<B��s���^�M��gi��j 9�������҈*��oD!jxLd7�h�}8�|ޞd�G�(yo��9�l�ٸ$ݫ|���!1Й��I_	`�ūX�"�T�hZ�]t�fx��#�K�������`��U*�ME��>,R���aP�Q� s�Z�Al�P!H#5����j�*��!�"F�L"2÷�	������[�������޿��sεo���,w?H9/^�a8��x�fm��}�.��J��ߧ�5�d�ڷUy�Ⱥ�0�ځ��.v򣣣�٢`cĈ��]����{��N�/˃���+����N]�w�;�
e2�۱]II)B�v"�d���Wɴ���E�y��JX�x~�2��n40$�J?Ȣ��&>W�xl6���,K������_�$&%��W�4������8{�t���@���ym۽���/?)
��럵��T�_�<�d2�@�ħ�*M,��h�q�̈'�>ߒ�-�p�&lK��폸�I !���2/�u���V��S�����_�ۮ�V\R2o�TpP\^�����A�?�ltp�־���zW]&�@rE������D<��8��6-�%O ��0����[����By��@�<��s� �Ո�L)�Π�����|ЙA��	y���`�Y�-�_�<��7>��x��7�h<X>��I��e�2*�v��V��Jv>:�序P|��ˣ�.����M
�\&�UB'U~��oT�/[�tϓ.�C����|��T��`�����y{���B��h�'�N��\�f��ۢ)���]4F���]�qv�;�Ν1؛ׯT�0<��K�7���R8y�+$�uO�����腚���jY��@��]A5g��@�UcZ=�ؙjd��hxm�� ��W?R���I�0�S�5���F~�}�*_Yf��L���W�����>�F������+V�)�%��Krf��.~���#y}��N�:�E�K�X!�o��Hkܼ�z�Fғ��߄�9���>��zwlӹ/lW l�N�a0<�xh�f5�}L1;xkY��<NFG�t�Z����s��}���w��M�0�f�ɜ�0�8O.Ȼ�y���������ߘ�xϺ��孻FFF����|�2�`�)�`��[�PϜǕ�9�Kw�Mb=�GQ�G�1���*�TN��I�rURa�щ�gt���ڪؑ�)xz����[YU5¤�]��O��W>Ag�I��~�.�����2A�I����<00 (d�k�dP �9�*N�:���$`�C�Z%o Amu4k�VU����ŀ�3ʽ�_k�<��bY��GGL�g�]���Vw**f���X�Ó�'>��֦����7@0�D)��>���ZXX�j�ÆWY�]h�x5�>=;���AǺ+;cG>5���E\��a���w�Qr�p��\�s�u��ѵ�ׇ��U!��c�Ox� -;��6�~��;��+���o޼�?>>>�����rӉ6&�\�J�p�8�;-�Ǎ��/�1`�@�x��&�_]�w�ch�����(�oQSS�z?����c�[o�2ue�� �z � 4*�Z���t?�|�qoPಟ �[��IXw��;��܃�S�����ܪ3T��7N��i��k�6e�U���H�5��� {(��\>��bW�.��hO�U:+8��\2���9�n�PWIee�Y�Թ�Nw^�����@X��lu���t�p#�!�2�����(��ȿk�J�����9�$)�[����p/I��c��ٹB��H������79��x��&$��Y����]�qv�xOϰM$�GK�����o�r��n��R˄/�T�u�(���Rxl��]P�dY�z4�MHѮ�4y��	��+5�e9U��:���{Co���$����B�C6�%<��s�஧���˧zF&���$(lɘ�ק@_2���#�;�-qT�F<�+u��5c���!,�W\�~���I�:m' �/{��$f���F`�@���O��mc�����)3!n�:[0w=C~3�j����Y]Z��3�
z��ձ�����.<�������w@���-Yz�{��`�kcB	�� �T�Hk��Z������2�������O"��C@k���ܔ���sލȧ��0f���y��j��T�����5�k�u,�1}�SQ��f1D$uǾ�� Cm_����HNNNy7�J��D�%ݥ�?{���
��� ���Ay]�^����3���r�P��V);w4��ݒ��.��p�Pk{�UYVZzV�݃,o4�=�j XiL��H�m�B��׺�~}�FkFo��Z�Ж�	�?�S�5���'���wSw��ͭtX�9%��l\�ٛ��"+g6�O����2Q��
�~*\a�I'�5"�d������O��U�����)`l�/�+��8ŞT���Z�́	�?N���A�~�R��
Pvっ����q��y�}�?�R"GEA8��C�C-q����.������ʈ,|�NO%xɻ��p5�k�Ÿ]��+���Ԛ
��q�#Ną��8��J��p�N��^�y+2픡�Ri��S�CxO���c $
ۘ�i�7�Y;q\���yFS3�WE�.pK&/���:��^�,�\��lܮs?fu��� �Ԉ�\&�B1��^��a�0^:���;;�8Ac���0U�z�j	`,�m'�W0u&0� W6X�
b�K�������
��'�$�nm`I����W��U�P ��˄��0],	��K����ޥYd:�5
S�^+�W��H���]<��:���S��x��F�����r�Z��p.�Ķ� ��ȈQ�צ��n����B�{�6�����X�@�3 yR���Kf��XIWxCW��" ��NHagO���P�E\n20�%.w��Q �=ť�� ֑iހ�22�j�A��(�K4��^O)��w8��][Z�w��5K�������^�+Q9y�'���������!d4k�j>b�!688���N��;��.ƣ��ʀ��]�z�,ʉ'�v��7Y}tg��~�3k43�q��F1�m��<�D�R�&_ʊ�Z؎/�X@��܌�|�;�`�U�N~#̮D6l�y_����
: x��g����E�k�/��ѫ� �i#IJ�g�t���Q-�|4����ҝݴŬ��,��lL!lT'�;:f� ��A%�6&�G-/��];�G �l��LCD
		麨����S�W����8�pX^��/��H�Ed��{�A��������k;��	�Jգ��Kh����Z�3j�
)�@����a)�(�\0��\�氞m�S�6�3���q�r�A*����.�r�q��D�&�� ҄�i2���O�,/lo9(o���<���+�#�D�� p��<`�+w�}r5�eq�S:�<�*��l|� ��o���Q<d��T������������{���"<�j�/o6RĲ$�V�i������V��h���`��9i�	�fKQ���Ƨ��2���077'��[�w��;�K�hV��

�����`��q�5}�y�v&�LfB�>����{Y��mɺC�b��2�����m@�E�{��u|�/c��4@�ં�'3-Y6�5��*(�8 W3 -O\��Z���	4]<;z��g��BI|�m�B ��r�3�o+���Hmm� �fڟ��5N#p󼩗J
��	
�1����|��?�����v8�P��*��{[�@(��8T����A|�M�������@	/"�ޘ{�BK��2}%1%���?��Ɍߕ!����F���y9>�
ɓ$������-,�� ��N�-����K�Z�!�p4�OEiH?{hq���
s�3X��Z�F�9�6;;� U��9~؂�a�3J��o�*��ۺ��b����0M�z�e��5P�m�I�œ,(�Ҳ�(�m�g�z�j��!�bV.`0<��rI�)���\T8)��
R�Ѹ;%���x3 g�x�r_��o埫�Í94�Q*���:�4�*���p�zO�);�zf�s�<�d���8�s���pxA�Oim���徂!��f�d3���Q	�?�w�f����Ə(� �/j��ʠc�!����K�/��3��^����s&����{+Wd ��̌��r&��gg�=����Mۇ�5�������@bo�ڷhhi+�.�(W�n�8w���� ��}f6�P����v�o��i	0����	��h��>�w��QJC�Q�- S�L}F�ȨQ�4N�gQA'W����|��ԽU�DeI�N�1������0DC�^0r�������I������g�52Q�mdʰ:�g� {mp�̒l�rS�m��e0��ٷ����l�j����7��w�ꉋ1HKXn��F&M�+�w��)�ş|���W}��ƺ���=�ɝ�T)��ow���X��|�s?/�A\�W5���� 1`���`�w�8t�a���RuO/?�u�4��׬���.Աpu���x���'ʐF3;lR���ɷ�~�m�����#���% l��7��:^wl߃��`dq�4��������r5�ߙ��F@��$�8����[%u� �O�M��r�U�#з�?7\�/�ٛ&Ä�B���J�8�lfY���١;8o�ܦP��?ّ X��fZ�2-�Z��C�S23h�����Zd�yǽbO!d�NZcԗut~�u�\��*v��f���,�ikM��JY�zi�U+p��O��1h�j�@����t� ��-"�=��8��e�����`�[�=
�%%&Wȍ��o)�`E������p�F�k�����������澒�bD�6]���4W��;*G�vBD�l,ٛe��/ٗ�����	Q��J��R�@�f劎@b5c���@7g ���U���uZ�2��2G��Z���ۋ�gkCr�&x�ůpD�S���*�eP�{�;�i�R��N�8����39�� 6w��T[�X�<���h@t�U�-D�6��ig����� cm��[��h%�Y�����PU`PЄ�e9(g�`ߥ��:(S�y��U�nԦ��]%��˛X�i�����սC�����:�U#�2�j����L=�oMߨ涁�!ո]Ȥ���	�P�W��+��o,7�ڐ�M����UtU��`��%n˸ZŔ�X����+%��Cr��@+�+.�'����ٙJ�G�����
=��uK^�f��]m�֝dXi��1���o�L�k��ɿ� �b�o�B�}T�}�:T͞7cmUW,�8P�e�� �5�kL���R=:]}�¯#S7���=��3��kS�l�y_ ��� � �RM�@��d��$@�VU��i��,Q���8cy�wo�$xI`�n��AFe���F�"������k�_�㌙�]i_s���V�;��B�}���O@���������f��{|���#�����K��@dzP�eP��A��WY�� ��5M��HW�뿧�D� S5.8�{�|�/,�Gv��FL������s�$��.��Oච��˨�im|L��O��6S9�elA"�]曃c�8����u��8[����X��k[�q�@@h�\&c�9��T�d�.��OJ�.�5(G����\��Ayǳ`rpa
X����񨑾�6�(�ց�4�䷟�Lf�o�Kt�M-U�9�?��ywЦJ��B�W���ȭ)��n,��o��;��a�jJ��������]e�J��N�?�a:������0Nõ[��iH'q�����R�%�2d�6����L&D��ލ�.�ut6q>^ؓ�EO"�#˛�V�e�����,��8��3��L��o�3�޽{�����͠�KQ�X�1�X�t�����?����S�G���T1�/e��u�-a(k�[5����nH&o�5kB7���L�,�ލ+�B�?:��zyz���&���b�>��>����
 Vv�r��*�����cu�rn6�7��R��N���������8���>+�)1^���3������R�,N��df���X�{�R��hз%8?��k�;qa&(O���@ؕɖ��p_�K���ˠ�e��'��!�.P� ���U_�-�����TdzB��.�I���d�ŀC�R���@x%���k���M����N89�U�iD��C�X�s۰��X"��@�pޠ�����v)dq}�~�X3Z4�f?����������EZ�W�[�ٷU���=(�{]��Ş
tn��101A:��t1ʍ��7.��):Gܱ��\�^d�	0S�=��^�&�9���[�Vp�\ɸ$�P�mg�p�^X�<ܣ+v H�J��rGg=�����Iw���2�z�����K���n���ۮ]�N�?_�]U��Ot�SY�]�d�C�������@�q���������Z6���<t�'�����T�8բN���,(U����O��@`r�Qx��<\(˕.���B�[nL�$�Ȉ,�MY�)_�mh�P���x@�8��dq)o�ӛx��4y?`|0��|�#�=Y\�~���ӛ��)�M��/풦1v�1�˕��t���]��1�䷒DD(Q9��U-�Z����r7��FU8�2bG�4]0���0�W�}��wO>A�gZ�P^�!�L��ч�3p���z��9vz�ja�Xb�,?PJ
+3um�F�bT�G��>�����%r��� �پ�Rqy�t�fm�ї��	���咹6��%`���1m;�-E�M�ݎ��<�h�x*�݄���b�J�H���3���=��%���zkd� �!�ʤv��=�q2�z_�%��UŌ�Jl��s�kI�tS���b|]<�M�~Z���k�!�ם?	:p����U8ܩ'W77�B�q봣Tq�eb<������,��T#�P�>�|��B�,y��%��?BD�A�׃�,:�W��-琐ܔ��iz��C����O���(���t Um�R C�S��	�3��,�_Z���t`�{���2�/^%!�2��U��j0��������,l��s�~j�R�qQQQ�(ϻ��w�C��s,Z��C�Cn�o�t6�	��K��`׊�����SG����}�s6�&hGr�� ]ɽ/�E�F��%0�� �D>���4#�E�;����8ם>Y2GF�b�����S�*,�w�u�mh�i�4"p�����@O�h���%���Ρ �1Z��[Y���Rh" A/iނ��X�0<��w+�2S���;�.?��wp�����-����@:�w>�����N�j��8�sN�g7��*���D�w�f�&3ە��ϖt�]"x�m����nC�}������l�|�WI9���,,��]�_;{��E���`��t���Q����P�<B"K===�k�́H!�/�(���.>Y}�Ӄgqu�N���:�e�y���7t �=��S/4
��ɏ��݆�W�ooJ�TV�� ���7H�q|���д�g;�`�A߆A��pBLg6��g�Yk E�@�SH6>��q��r6B�;��#(�{�\�KȚ��8=����A	��AH�@����qi��9u1�lrP��<AU���[�S �Mf�nk� ��Ni�~��K��?�߽y:a
]s��MV�d��$r�O'Iz��t���M�
�V���$J��lc�]<����5 ����?	϶ѥ���Ubo3.7~JzN\� d_�S5�b3N�/�� ��O��&|�Ɩ_<ZQQ�-�oA�g����᪢��|�FEH���R\��F�l��� �,G���p�# 7
������@���3�/q~�,�w����tj�q��_	�����괞�'B�7�9��Q �e�O��D;��\�1�	�T�C��r��m��E(9*U  �	>1�KF��d�@c���
�=faȷ�{f�]�0222.##s�&������$�IBI>*�R �U7YOrrrpi���� �q�;��B�9&�r~�LZ}��;#w�R]�w���u�L�?ԅs,�V���j������Y�^	J$�7+�	IF��=�ܝ��a��P�q6Ó?����J\��M�kp�%����ʸ����N�j&*���>�;/����a*�ol;?�a=�*�(��C%��o�wvιj֞�΀��	��=48vǖ���~T��Ķ�d����Z��>��Z��'?���/Nz�[�_6g��<+T%�s���h�p*��ȚX�sS��z��{�<���������w�w���ocj�J<�22:����︿�|~Dh�L��D��:Ď�Q���ju=�w- ��� :=H���c݇Ǧg��d֗�� ����:ئ.Z�CY ������9e��Ci���h��w=˓,_��7�{h�1�^7X�+R���-��?-a�6�TG?�Q:ՈɆ�������� ��d� фd��Չ�*w0�O�=�z�v�pt���gȯ�Km���U(;q2�����pk����W�;.h ��%����ꁣ�hu�����%�?�
���C3�DљNU�άt��-�e�gJ�2�?R�n�G������cg{�Z�bB@=�< h/��I���W��s�?�Ǘ�>�/���tu'Z���=YѺ�{5g'N|�q����8nI�d*eG���@�_�Qe���0O�����%@�p!�0厫j�2�!�v�w�_
��ne����fm3���fm����v�͘ni&#�,$M���m��I��)DK8��T�eԬ�
/�ؓ�a���De�8���u܍S�)���l u��y��N7ʒ��~JF	᭓d��Pۘ�96<�g����{i7D����x�2�D��j�S�rT1j��o�� �@�_,��i�i EdE?}��_-�ޠ�4)k=�)~�V��H���#��g�k�?	�1]|�U��~*��2k�~Q�M�]��г6���m�|���d(�,g��o���F�s=c㹣�ć|���͆����������o	-L�-��&�����ޝ�N�>�#�j���/i��u�����ݽ�\�;t���*��'�"IJ�����櫛m��b���?Nφ��%�*h1�U��b�����z���@͓֙{�:7W��w�E�H��O̗ũ�2�^e r5@���4|ZIy���|�rʕ�YLd���ލi_�;QmsJ?5����Î+�=��D�؎ѲkP���k�����3�i�.�ZE�(	ᓪ��!W�>y���{������ �>�	���H`g�S��ե(��sVo�ݾ�ŠJg�$@t<	S��vJ��G�Oij�/��Um�/ ���|1�U����u��g�S����o{7j<c�xͽ���e�L	��,D�.�D�y�p_����d��=Mޠ�೎��V�N��U�^4�P���rgձ���3Փ��^*-�*�!ֈg|}}9���N��s�G z���K���Āv�Ş�R~d�
����7s�C&dI�+�6B�� q�1�A�P�1P�}��V�]��b#]=��_ɳ���7LܱՁ&_�X�i��p� @����T���ů��Θ�<i7m��2-ŵ.��}�o)���������P�!�q'�3&��'��=(�/�RS��!Y���'MxJ3��}is�y�S
15&U�s��1��W������ų��^�-^'�s��~�0�Ŋ=���g��Ņ������x(Z�Oe��A1�{��eJ�h�;?�6.�'o$u=����!�?P���y�T�vtR6��oHk�yc�cPu����38sAO�=������-�}x�V'٬��ص�ؼ��-V��'0H5�Vi��咑�������y�u�6��\������Ş���'a|��58r~%��{���av�ǜ�)�.D�u�>ٜ�~ك>���F��L�5�6�������VVQ�$���V��sظ�����#�=�ʂu��gPpt)�-$uWR9��%%�ѯɔ`�]ŵ�^_з+����U0U��ԃ��[G�V:��׷Lp6Ğ��W������_z2+�,"ˌ�y�Z���U\@�| >�h2^��Y=���2g���;��k?�0���KU4��m�֝��]S	8��s|P2��;�!h���j�J:񋣠�*"��4�­x��g�X���ԩF Ow�s�2(�OQy��϶i5`�=����[��$&�Y�J��xo��ܐP�+5����/�7N�q�-m���
h�1�yC�B�| �b��kQ��+�r����ut���N5cH��+�g�ݻw����Z��a�	��ac�J�~�m�	t8y��3�(�����V;"o�fo;Y�L�`�J~;���[}�/_�\l���ř���À?~��Bօw�r��+���#K�,�W�ݻ0ݾ?(�]9����K�ζ��T�
, ��c��*��U��OS�+�FA�e�Vra���D��}��]1bV�x�`rj�T����L	���-��/?*���P.8�����u���Б�Y���ok1�'M�W�� 7�0
C�*(�8����7V��$�ʡJ�hr�X.����2}�eyy��G���r�e���1�6p~S}�@Oo�`	?��-9*��p}&�/c��N�@s���uO��X���4���1�s���}��$�(�/���2��Y���n*���{_P�_~��PP1�mf6B�y/�s�ؓ	�U�9~����'��ekJ�=����P�(�͏<e+y
8c+��R�nC������������L�_����|/��C�;��C�`�N
{���Ϻk�T4I��Rp��ڮL��X���"�Z�[Z[[M�P�$�,� �4������e�O	���)�V�C㝪�� ���wh��2��'ෆ;�,�Ğ|X���	�Ne��l?MN��~:`�R@s�բ��w}I�dsX����
��$����%C��JFMM-r��rS�'\o{F5H�Sr}S�k�����y�~W�ůs�� tl�>?w�
	���6(�~���Q^���!9�-r�W��3�޺����ҶJ+Fr-��%�����zÍ�D}��bG���Y��Ќ|b���MB@�#������o?V����nB�����,����ۗ�<�+ w�at[�Z���#	�����"���H�q�&S�m´
�B�{$�ᤷʚ53P�v��K�Ge�%AF�v�a[J�q�e?`����N����5��r��O��=���}Ͼu���H_|f�C/,�6<�\���F����Ľ�#�0��,d5(EhE
��7`�8 �5����I��m;��Rt�)�A�^�'�QL��%jTM�g�#�G���/� ��`& �(�U�ʔ�&T��q�.�����o0�^���_�l$��K��tHS~��zt�S��p�]".��	[�/��g���b~-cu(��=I[�>�.�v6Ny�f9�3(���`,�cR�ke/���������N��*���<D��>oL�X����*u�N~�	�cJ�� d��||���
#��iX`�sp��rT�$/��&��v��V�	�%�&Ը�~ɄD�%O8�_?�z�S!i��y�w���uLI�9N4.7E7mB�B�;_�t�9�V�eq��(�y�}C����9a���)\��l�#{�����+?�7�+��V��Y���-���y������x0�q|�vO�F˨j����;�(Ʋs�Z����w1��`1��[�b���Ѻ����LO�r|�����h3�P�ᜈ8�i�%��/qk���R�V5�I�b�+�2l:n�q�������NB1f�hY��.��/aϑ�W����tu�xP~m�̊��F�d��n�>\(�[ڮ&��ҷ?R�Vk�j(�2��6w��Wސh�/>a� �S����i<�ߟ|"�α��S����|n#<g��h� �:�:�yh�!f��z�-=C}��WP�����m��T�՟Q�-�;�僝~���>��Z����<Yh��T�]�������6��t����۬g+����o�p�XP>���Ѭ�@;<��zr�m.G=z^�K��ϙP;{����$wg�����6������qx	�.G��.}��=��`c�e�ZL�O��ܓR?�.w�@"��Qh����Q���Í��Yw���gKAt��6��
J�2W4ڤLIy�hÇ>v�N>�B>�7p�u�2p���&<���0N/sX�8�dl�!��A�-`��8%���x���/�!�h��ˌV�f�y5��c���``ǀ�C�c=��_^.~(���6�>	PB�"\�X�5�;������p�e��r9t�_^���t7n�e�B�#��Q��3 �q��$��t�����I�ʻ؁�.q��~��3rJkj���;����O
BkVA{ד?3�~T�m[�db�6��U�'�����a]-d8�Âkf�G�d+$V�Q�����Af@�D4��j�(cH��,�}e��?00y.�˳�'SÏdU�P�V	$����� Yx� /n���|[|�a��ɣ�h���%i1����#9�����ɇcwe���)��wݜ�)�{4�&�h�	�fd)m�K���7�p}���ۘE�5�Dk�ӝ{gF�6�{k�S$�����s��_��\�KI�D�R�<cW%��!"��ѷ����C�kM��׬aǐ�D���#�}5�<RG��_t8�������#�lqPN�|Fw-�Wz�t����8L��{�����i��w2����kTT�#�S;/�/`�J�؅?��W j�]:��LZ}[����X���f(l�,y&JK��N%ߺD�V^O�5��^o�6o�+�<y
�0��ַ�ɫ�J��:�x�*+҅�7י�]�~۽��{��ʎ���M��sZNWt��u_�oc¼�R��;���M��e����51]/���B���xX>�oЌ��]\�����I�.��Z��p���Ɍ+~sB���[�ZS�`��g��'�23�.�W�	�L�:��8���x�UA�-���
��
�V�����T��\��O�g���^��U��.�e���xT3{Ԑ��c�M֜�}�ip�W1Z{4�G{���2�����-���,u��A#�2�3}f�ۇ�n=���q�i���b#��B*��Oݱ�4)��vKjY���j��qħl��`*'�W�)>��w��=H��VO���}&d���v,�Y�j��+g�T�/��=!`���m"�g^%���j*g�Gw�1�o(]����R�<)|��J�Ξ�涣k7�����(mrK~�Uq�Q?uМ����
��*��E��9E��!���'���gv�1cP���6����g��v�u���~�l��DH���e�[� ��pٟ�'&&\A���	��7��}yyU�!Ls�&?�0#=$$wh��S_����p� q�� ���oU�OG��}�eh|^ac���%h������]�Ǧg��w�B.��yА�3���,����C���26@1i X���]�:�����s«� L��!	i�W@+��l����aj�q��\OX����mr�q5F��@�ە� #u�$&�/q�Є3:�A���a�I��`%��"�����uLk*�qSSJL/��x�xͧ�F�i_2@�]9��^h����p����#��E��F��&��Mw�!�X�;(�֨&�x�Vq�+R(�U������Kd@d�=�ŉ�����MC���q�e�n��z��� C�x��ލU�2QCfx�e�Ɨ׵9��,֌u�9-�:k,�i�rps}\n1$R�S̈}D7D��@����kq%�y�㬞��Ծm�X�pH�;O��L���p�T L/hcV#	�ߧ�*m�̾H|��@�N�ʧ�����hp�9$�KL��%���F�*��L0X`� |o+_��16GMOxV<"%� �t [2�x���_��!:'''��Y�
P�mg]aT�qX(H)�����^������{Q�o��2)x's��u/:<0J�IK%>Bs�L�%2��7�!��6	~���?��r�,+!�x��ZN�W1���L�B�kx����nX�U|
~�]�P�Љ��F(O�k�)�`�؛��j�l�K~����D��A�x3f�]���R6v�r�VC��vm1�u��-��^ �;���,���\l``��`�iwq[Z���R�$	I(�@˃CCC? $�9����+ݠ;�Kh�I�V��!1I�e��x,�}y�Z]��Ɛږ;駆�p��w� 	Mq���aE����w��ҨG�Xb̤djp>
�~ʨ�N���~Z1�6e��f�ޱ4�y����{���*�LC7Yb,�5�#Xo&H���븰D���h'`q�%8����2��l+9##�Y�]�6���u�@��/�En�A:T��Ʒ�p!Ȣ��ܢl�j!���ե\���8b��ea���E�m��R��$\o����_���� ��7�YI�J�N��$�W��M4-�iSp=�˅��n
�	rKQ��y�z��j�����f�/��r@�f��.�'HrF\){2��uŢd؁��sؽĒ��NFwf�|e���z�xЌ'�K$��B�����>����WJ�~h��i�c-
���I�5gެU(N��������
W����g�K��B_U�]���F��ש>��4�g��b���]¬�Ĭ��h���~�DI �� ��p�S�Hh�;|y���禯�JR�9$4i�\�!�\�x?>�hnNa�{|�Xo������r���O��B(>UK�qH�&���a���52>z�gr�I2H����k	�ח��+x d:����	������
�,K:_�r��L�-x2�Zz��O)�r�AX�&�;���X/�]@��!���Ր�*
4�X��������L�P:�pr ��䰦|qf���ъ�\.���gC�i`\ L>���K��p��:�/�D	�Ĝj�)���ˑ����������ɧT�׫����f6&c��+W�nC�@F�<ÏE@�-�vV�wNӑ.���_�Vg��l���X�KĊ�"��@�g��'���x���^�&	k�c�U�Zcϐ1��N8�׃���	�Y5/&s܉���Gm�/�ˁO`,"���w7��Trm�7�1��m^%FO8��7�1+U}i���Py���T��ɜ&C'K����>)�3��毟�P�a�}�U��R��H��;�?��C�0��x0�hO>&AY�q[�--E������ޥSm����f}���?~� �dn���K�9�������P��/Ep!��2�� ��PQc�Ayn�����L C�{�ӫ�n�:�O� )ܳ*l��p��R({7�	��Ҭ�������ȅ���?1t����8 [�5����w b���N���e����ٝU��
����~oeL�k 䌒h�i�]G';�����{��7l#�xJ�B�e��f-���kA���pN+�J'f��4���C�! #��"�D���ma�:Uy�Թ��zb����p�A0v�v�3ڂLVh�PWBx���MKq�\�[����=���s����^�皤e"�?��j��TꜪ�|��+��G������_CZ�Wgg�J����1 ]C&��O��G���bj��p� �9�/��OB��AHƽ���L;�=��z��˗/��ÕjZG�wɱ����h�qx;�K���A0�ղ8��L�[�fOO�Nfs_ܻ�D
���-���X�_=���@ZX�-�[�%��؜� Cc�Ȉ�l��t"���r�v�K��q���duN�Efյ�m����V��JjQ(J���H����!����O2���zUzD3��XQ&*�"�lR��UK_�/(���� ��X�aط�YG�K[ׅw��O�,�"� �E���䊧DI��bE�3�����7�7Y!� g�oS�z�"���#u�����J����f"����`3�zK[�&I�Lk�J2BQ�ۀ�Y�����,��s?��o;28������aH�4�}����Kh�jE�Jc+cZx=FH�����Bb/wat�zӏ����d��L���8Ѕ�z}�X���͇�.(�� W�y��q��`T�lY�����
�IԒo�3�a�0�����{��S��V�_Ǳ9�/��,B��v�6�2��x�MBy׷=�����	؄2�	!Sw͜1N����܄_,ÎU?>��4��`dsAE.�L�N���O�)��O�%=��=k�9%_r�哂�e��;��,x����,)sss�Uf�d����jU�UF��`@�����]�f����6���5�y#� �����+)�Rnܩ�����\���*�mS98���8�������dA��󤍡[��ҽ�
H�Lww�)�C@q8��(��d!�r�f��]{,�PN�M�q�_%���>}�̘�'M�>�!��D`c��q�i{��vG f~��
���	!|:ʄ�){�\ f��h&i��D�$"�N&�k(�*5�eI�A��m%�&Z�oƷ��/Q������3Y��kZ`��a�hY�����ǩ�%���m`�u��G�:;�x��hl]���f��ꂡ�����B�\v��|���9�m
 s���aLC�!l$n�Z�k ����j�2��b��3��	�ߕ{\��T�WA����Q�g>�.�=�Oa�\@;�j!�HS�h	V����'��%=�xn���4�,ib�@ �M^�[�}�˽�J��8�]��������	 ڀR����_��$+����U�ɤ^O��
O�Xx"=�ֈ�%r�[�M��j��ZB���r� R���61�:��a7:���D� oS"�˦G�}����%��'�؆�fUgF�m�y
��K~���X���+B�2�IW�f=�
���F<��H�6~��E[�|&���p�+�9��h�]p�?�C����[+.�	C�@�nA��Kr*VIǫ�$F���vK%>�ןΩ�1��?�kM������9I�t�������/� �i0�cF���[g��� �_�x����Hֳ7`Q]��YH?=�t�C՜��}UA��Ц�N�Hw������I��9��N.������X��u�Ƃ5n��`��&-��<����+��\�G��
E$�c.�e��㋚������w2���QQF�;_�:��b=ۉp$nB�n���bI�$�-޿K�����L|�N�'(֚���v�������V?�5��(Uժv���b�Ӯރ�ܡ'��B�{*i�jR4���+$r+�?@���N��������\���A�r�;=� ���hZ�-���&"Vz�����腓&���(�M�n`�\.@@d�2yYԣ��c�־��
e3���+R /~sl:��VȲ�}�{����rv�D�ba?��9����c�I���!�^�m������Y�}�~����	�4�Y�(�#�Q�1��!gvp���閌���'�m�RsMJ<I��}v�HJ4x�!�c�:.�?/��tLమ���?�_8��c�n��:�!����lNg��y�Q!Ό�#�����%��4�ϯ �V6-�~��g��FJī�j!bxօca���P�`���l��>{PNO�3��DBMc '_�d� ��8��?b҃������&���ύ뙋1���?����GD"��C�J�!jhy���b��{h�o�Yb2H�U%������Q�y�Q��p�+2�hl��Y�9������ݨV�0�pF�ǝ<� ��#�m)�0{䝔��v��4![A\���z�6���	��/��N5"�zt*\HM�p-o9-��\������ ΅	_=W�40���RɍB�7w�A`�t���JQZ��҇X؋S`��0��ӆE��/ɐ~���o� �eF�r�ɿ��k�ZhX[�l?N�b�	5Z��v��?@��*9�h���(�x��(81u_ !+º���J�h�����7Y� ���H�Q��J�$��^�=*�����\�W�  �몞�cy"� oP���W.�Pq��i���P09 ��v��$|�ގNJ��HҨ{T��~��"�f�I��Z��p��ć�M��x3s�H�����?5$�0ݟ�1�_�x�3���lh\��4�
었=j���0*'s��j��v���C���a_h�t1Tq�wzp/�t�U����X_6�2��r���o�C� ��>]���9�Ӓ��R"��Ȅ��E����HJ^��v=R��@��<�m�Қʻ��v!%��g�����%[/|��s���>��Jv�dh�ε���ĵ��&��'�?Qhz8*�|^�Gk �XHE0��E�BQ���?j��^%�D��|��}�_����Wټ'�W��5�y�䓫����o�-���p���_?�<� r�E���)�`q`u���1�8�PM�lG��H�C0��J��
@#�^v(P��"�����t��.C�b0\٥���{�^x�E樭�d~%$�*ʆ�1�o8�����	�待�FB������(��Lֳ���̅��eq���3��=*~
{��i��
 �I.74J¢�Ķ�}��*]�d�	9Iǂ1s"]�,��ג�Ǽ�J�2P�4�:h���o-4�־ѽ��i���1Z&d�7�;���.�=nZ�g7q��]U��F%!K��na
�ؖ���4p5Q��bΣ��e��χǱJZ"�s�.�"M�C����P%�k�xy������i�:򐢒�&�y�`��m,0��mM���o�-��b�5zZ�/H�ns��A�%������P�*c|?#N�3��G1=��Ȑpi{�l�c#���dRȝm���<���$��cmwUN{�CA{���U�X�wcB��|�A14�˭����Fp*$d�1�r3^��<�������gDu��WH,�}��]��}u>.�Y,��������s��fa�b������@�s\�>��ԩ�[�~_�A�q������4���jf�H3��[��"gY�K�ƟH�u��K��%�"�Kv@`���"뉜��R-2��yD&wSUd�Wd�,}���j�W�j6�N͎���G��8���5�x";�� }#<Z|8g6�L��{��ލId�^ͻO
hi8i߽���_�a�Ɯ�psf:�[�+2�4v�29�����m�։�V8a4�{&�W_k�7שN=]e0Z��Z�F���vR���O���y�����JB��$le�5��x%�P�����z�\��G���U"r��;�{@�����((�@\�Ap�v�&@
W�o������^�Z-����1i 5�����)CՅ�fm�|��%qr�c�]�Ľ����YtZ���<Т����� �@�:�T@����U�D��L�u��6ߞ&o�Љӏ��`>��HP�'�R�L�4����cp�tt���-��tP�1�8��ri�V�ҥt�'�q2�#�?0�
���B�I�= !='�]����{�r|<Y��_�蹦l�D~o+Aɖ�dZ�E\.X���'�U�o][`����w�*8/��>`�a�w��vj�ec:K;nO����O�^��%��	�g��΀���d��:�0����2��Pk�]��X/{4x�צ�]��й�\��W?�� �W�bvp�_zI�";kv��6�C� �B�������p(g�F��h���/��J�U1�����J��h�- ��[Λ�P(��Z����s�r���;r-2�-���	����t6ΞE�%Qyڻ�:**�G����	�����dm�e�ÿE�C���|>`��s�[��/3�輾PGEw���[��q�uutpO�N?H�]���E�S����ɖt��ыc�ٔm��)ؖUc3��OI������y<U��~��B�R�LE�S�DQ)���Ǎ�*$��
ɔ�c	J汤c<�y�=k�sNw������{�>����Y{���������{��诎,�jLU��	>O��͝D�B�}�}L�У��H�O��K�z�Xl�~���K�����؆O�M�R����.h"�~��+�t�H 
��#��?\1gH�B��
�v�	��8�V����T����.+D��W�v�H���]S������q�����A�e�4����؂�OH@�����ja��\Օ���>��D�f�s��e��9
��H�fS���x�I�(K�c��S)#��(c��3<�RP�t;d�ݦw�~Zm��p��P�L�V���c�!v�>������k2؅�y@!c�ߟ�ֻM*J�!���k>]?xG�$K����A�cZ+�A7��`��@bO4U ��|�^\�h�ƕ�I���un���q>G��##죜e.��~���q�uGvb�_�J����������X�腤#q�R�<==��� �	|��\8?�(Sr�Uׅ���C�g��{Ze���&�Un��>��eР#p݇1F��Z1�"i��)�p+ܚ�6�vni�kE}#P�X�BS'\ʶ
<��gP���Y�m���P�\�l-)7��{nB��j0	�����W7�d��\P�.""R�� C��{|��nT�M���l�ٽڢ���I'�Y	
���i�h^�ؑ酥Jߋ
y5FZ��Np_���8u���t�5�&"��*#�\jv0l�ĮU�kw[3�H���s=��Tm<a=�QQAS���ǋ��Qh��|X�߬���������U�ݕy��f�xC	>��؇hL��j9֐�n>� V&��!9����5׿�){g�&�dV29���X�^�����V[,�{��n)����X�)�U�5��t�ITo����m�[���s`J�&��F�z$�s��mj��::�v���Ô��nh{�f���[3�J�\�в�Ǐw�r������j�`�)�䉈��Hu�oE��Y&`�V��e+'Q�� ��a��xܟ�g]ݶ�\D=��y,/�-h������|���h��r��e?� YC�[�\�C�vb%���b�ׁR��N�w�$Wk��
�t��_�P:�u��� Uc�0�ᶰ�l�O��v�沾�5�P8�\{h@�Vq�F-�cbb"�, �k��
�ek�/��/Wc�tU����������kzǾK�LSZS���J�%�Ã�b��F��;���x�F�����Q����Bh���zbh�!�]������t�EH��E+	�[+����	�`C�t��D.g��Z.F�Q�8Z[��o�n�2�.�{/�A|��^�#ga�I��

�(�9���%�0V|{��T��z�D��_O�F�pd�ۑ$�ؠc�K��}�����@bJ�����\|e��]�����A�^�뼗"��1��������u�7�˿)�3�S��*�6jD��r�W�<�
���;c���=%Z�<���"qX_P$Ol(�M�>k�-�#ia�0��l���0F҄��%Rm�B��*Bw�f4�J&�i^�;�R��i�7+IU�a3<ʝ��"d�D�3h��&��±����M��s���ۀ)ڤ�9^��'�������e�=��76|b���*Ci����W�AO��=�߳��e�3,�vx;>�3���鼑g��G�?�}>|6@�1Ä0, ��J	n�M<���h��gAm��ryA�B\�0,!^�+��l��/!Hێ��<Ӭt�Xs�#�U�]�ᙅ
@u�T*z�a��8ĺ���Jx������f_����%Q�l_��M�,,u��f�bg�3���Sw,Pu��J2���Ų��?�b����M�a����d�\R6�+Gy��J��ZAsY`I�H�q�cn:�I<��|��w+�E]���<�~�8{?f�؇|^(��o�i�Q�����־[\��h���wg�ʥHi����7���9ԁ�[� ��Mc!1�{j9��!_��9;���,ļ�A�����(
�t/մ���ev!��b����ٝ�(:�iJ��o2��e ��c!z�l�]���V����R�æfH���IG��Dm[wY�	�H����EO놓�f(���l�-��v��,Um������C�4$}ꤌ�b�>���Ƃ��XO9��%���@�W!V���eQ��u^�4@g��1�@�a=C��``g¥l�MX�U�E��+k��:B>=
�����g�q�I�w���&$���X0�G$?�q�b�ޅ��i�-��28j�� ���$����| �́��5�Eb�(�:�}ؾ%����
Q65� �chF.�ŋ�oC���	r(��\��<ע��C���v<mE �j)�?�&��8H���	J�[�X��=i���P�]��w�0d�:��Lĕ�=������7�I?����
�Ny�s5ٮ*��AW���hP���2Ԓ�M#��T]�5WW
�^U���e
cn��F(�C��)�s�	h\ߧ�;�<�$;C�P�I�oͦ; �I�^>�|�᱇c���̡O;�
��Z/�h�����d]0q���G�G��L�)u�=YP ������[��{�g���z��X�]��$y�m��P�߭h���Y�U�t#z���f���e��;��\7�j��5�*�_M�(��[�$�T)g8k���*.��b6�"��^��:,�ZN���F�� $>���@q��5RK��gKw�@RC�/^����o2�������G��}M �J�� )��a�)��M�����ITfmD��I=������2����J���˳��}�ɶ��|�A]�t"U1��z���0��@���T�S����z=_{R�鱚�4�����;#�
�9A>�ѣ $���c��l!�O{����%0���-r�Pi��I���b� }���3q��!`��h��ᑑ�i��^�:�0�Զa��L��|��܄a�o��+�{0�;�E��b��$g<�w�S��e��L�L���:hՄ����M�ô)7vz��c��$LmZ)�2�F��|��,��SFn{9���(�A�{A�S<�.M;	�G0Y?;!�A�F��RKɁ}�ss92G	D3GVEA6�^���XIr��S,ĎH�����_�J�Q��ps`��u7��V
��u?�A��<�$���>���:�6�r��|II���b'g~'�0P�J�����p�����A�ډ	
��5U�E��gwm����Hܲ���mj�b�QzpF))�X��D��,$�xQ�>�/%u8O,�M��	}X"�}�����!]IHTE��I;��u_C�ڈ�{T �Vo�lC�X"[��Hq�K�jp����I�&d3C��I����z����1�޴�/5u�.�V�篠d5���4����{*��f`\-��̩}e��P,�Ӭ��jT99B�J���HC_sqNO�P�Px�=\T�����#�s�Ά	Yp+��S�L��J0V��H���q�,�����:@rn߼����+�[M}5Y�f�5�D3,���2��f/��Ր �>r�t ������BII��wP�� �Ky��E!�gx9(/�2�|�� �ěE�x�(�PN%�QN�:Μ�W!�,9�62C��,V�Qd
,�����_p�r�Iʯ�Z��#���|Oa��Ơcz��Ux[q�~9D�E�����*nSmc�c�ވbe�M�RJ�c`� ܨ@-�6��!a��M4�܄"�pC)`�� +\�#�{"��J��`��C1줪� %Y�w5>�"�s`��|F�Y=�`U�J�v��s��D�^�x�{�/��IQQ���s�9�"ŭ̥hBkV	�@�fv�w ���-b���WQo����:8Iυ^C�9i.��?!X������ÕJ�V>��HsqW9T(��:����.��%�0\��>�Ts>���6T3�hZEp�Wx:�x���cG$}��b<>:��GK��.񣾞�O�8��V�N��HJ�_�^����<)buސ�!p��Iw�3(����Y�B� JI�C�9M@Up鉭%[���e����Ao!I%��ډ7բ,"�>R;�I(�r��W�������s��)hIBVb�ɢl��#74����}�Y���D��jj���5��WcU�U��TT��9�p�MX����.Fj�P�}��l�����e����'PAck�H5F���8���舢U��O��Z���Pt7FM����q�M�R��}t/��6ˢ��M�b3���p)�xs�����t'Z�g��@l�(�hM߶���znL�b�麅�S��������#�2e�0i�L�&<*RW�����NM�UXq]��R<��ϔ���&�;>M�)h�K��c���Y+�8��Cl���.Q�`�xG��\F
f�4�]%7����L����˛��چ��N���UG kB�*������2���Xj�v|-���ީ�w>K�@��H|�2��1́o��Q����m?�s��nBxz�|��|��b理5k�a��[pSs�����#8�A�'7�t6�=Z/(����M`T����z�ގ$9B2$�Am����)o�ȱ%�a�ނ���M�%���1jU�.s�@��F�&�� ����1��|Jb=�0����A)Z8�
�k֨
�P�ƶ�"9Z�f��T��\�T ��0�M�be.V�R�.
��rz�%8A���C�WX�Z�WJ�P$Bqkv�	��5d��|BoB(�2��N!�HL̡*�����!{��H~�G�C?��pގ�,9��	_��V^M���n�8!���@��3��j N�t�`�'P>�TY�Pi�޲>�̈́�m�0�d��"yxA�44�YF�}7��wʺ��. ���~C6`��<
@b�.Y�W\�̡NFD��j��x��g+�zPF���	Q��ԙ�0�f�HS{%�\�E(VE(c�R�s�~(�\r�����+��O���9���T����Ji0X3����$i���@�"����GsHWX[�B5Zoۆ]7�\�$�Yyz�{to�������*	��x����"u�����C���aX�V���PMa��Bf�cᕷۉb(&|"��|� ;�cMD�ɵ��7���#5:ٚK!��1֨m�1�y�C�Л@E�/ �;���#M4��3�S�&dG�HM����qZ��{4��܃z||�w��Թ��z�I�Gb���o8�(��2q<L�s��c�����̫ E���"՘��^
�P	��赇ˇ������/��G��#v��ǃ/�o������xmZL�P�#��ky���3�j* ����ԃ��Tc���E��k�W|e}]k�E�e�4#�M�B*��H��O�Me E!��ԸXsg_l_� 2F�n"	��Jȫ�65>�ʀ�h����o�%��4�N~��ޢ:�n�h�P�����s���w ��WJQ�Ձ$��JGٌ���<��� �7�a͜������A��X=S�n� ��x��s��c��[�sC�ч���>����V%Si>(xΎ'^��*��(�ؾ�qtޤ���:���y��7A6�Gq�N�"�ɯYnή_�)�FC�6>k��U��+
��Zl|����U����ʐ#6��L ��Ύ��cZ�K���"i��ƍ���!��gkW�����M 1�^��n��m��z��V��56�mH��l�Y�w��6=�����Xߛ������-��y N�q�w:������X�P �v��#4Ҿϻ�k|^��S$��2��7(s�F�8?��d����A7P]T\E�-���g����2Hӆ:��5-��CS�B��W챬����צI=�u�s5!�����{�2�`��̲l��+�A4}�?+A�k��)d~�����v@��c�S�G����MWs���d���~_��eÁ����F0��kf�vr[�Ү'_��}u��������{ʴӐ����Ⱦ��k��?�X���
Y�KF�<2�Z#��u+����ւ;�m�����u����@��HSEČ@�.�و�\�?�3��h����н��U�?*e*�"�:/��,O�^M ��r�&�Q_�'n\{�O_b���bv7���#J5FHa����Ѱ�����Ԁ�&o�|�*���n=�܎�3�D	�G�������~�ߏ��~$�Tu(���8D�-�OmZ}ZcO��⺇t��8��"�OQM󋟌MU����h���X����]=zϘ���4~�?�u��ٛ{�����M<��hQ��%�U�Q��pt�ӾضsDj�#Ƶ�_�!��gb���+�*��wq�l�����]7���^���������]��K�?si�i��˧�������ePr�ˎ�X�KHNNVB�Y��W��P�h�0k����Ǩ�*�&JYu�F:�OՏN^W�T�bR���i�_F���C����U"�Ý.��o�R��o��,F��<59�>88�pN(��1���(��7�y�{ү����b/����ܻwϽ��C�;C<뺁��M9αƞ<y����´L����j�&����&���G]\\�ǀF[h�������0p�jp�t���je�Y���9���%E!jq����h?�H�Ύv�V�_<������纵k׺gx�,{��Nu�J�;R&����>n%-/�E��¯���P��w��o˼]u{������Jzzz7��f�n߾=�ۗ���o�98$M��uݾyS�z�ȯ�+�ʦ�~Qu�P��PTM�ի��z۬���c����n�9M�V~aȻ�[qʯ!����r�)����J��1�@�^��]����7�Z.�u������v����٠
���և�e�D���	=�{��y(+j&���ye�|���c�jWW��ٲ�h��jv�o�d�R�D�Z��!w,X`n3=I��膍����e^)���K����hR>���͝�����[�edh�)�`^�;�{���ܖei(c?�5�P�A���i����j9�p��h��4�7��$��������]>h��)��7���r��`����L*Ev���7b��e �ˮ??�u���c��0=��<J��kK�y���;Ff'��8���;��J>���/�n��u�K:�\%�T���V~�E��Ƥغ��n���aq�Q�量+1�"#���f�>�����
��m���s��Ϛ2�p���b��c��)������C���
��s�g���Mz�f�����v��H��)��8+�����#��Z����22.5���z"!�eee��UW��kփK3]�t_�"##=$�gc븽G�߇zzz�<S����S �'Qko�i�� ��o>+&	Z��v,{α��SVV��E7�<;;��B`��Q]f��t�;��������xw����2ه4�!�+�
�(���T�hh�<������	---3#]
[s�k����k��������Mj��#�@��`��촴���X1hD`�!�[�ܗ�Ә�EˆGM�K��ι��IۡX�*ܫ��iCGG��f�&�fv����˗/7�/��Ɏ�����>�k��]=Š`��p�ެ�'���'��+o2�[G�}�����L����{{�<��^���Xl�e��2ao��������G��E��JQHH���������p�J��ğ��K���t� P���'jZ�M<��|��m�7���&�QU��: ���Xؘni�u�Б#S�?~�������ӨE����8T4k�u�֒X��Pd�V@�d�-��hg]��Rs�Qy����G^���`����@���הEB\���e����=O8th"�"P�<�͡U��\�����S~���ﲲ,�Y�,uy�**ZQbbƈi��ĎvHF�����69�s��8�U�h�Y<".&6� � ӋLP��k���k7y����RXX(��³h�Ql4�mB��]�����d��ڙ�[2�۫��D;�<V�������9W�v�����.8:� �t%��WɹL�r`u �.!�p4x�l.��Fw�������J�9���W=:���/5�Bwz����`:ˑ�<G1;&?#��8 ��mxg8�~t+����L����Ǟ/����mg>s�l��x�<�Uo�os�C����C�l���)0��Ç�W���gQB�JQ=�G �M+,��6ض޻#F/����e��\歙 �u�� dT�#��7lX���#���oL�S=v��!�0��K�Di������|���煃U\�xLO6�ʰ�v�*��T,0J�n���=�W���i�egg'g�1S�<��K<\\���AXZU|��GEna6_�}ripp�iuu��>����ѡIo�=��������障�Q��#�%iu%7%ed�t\�5�SB��ϫ��.���c��Q�c���'�w���FejldddГ�\��B�YqF��c�������]_�%�<�O��HH�m���|���I�\���KGr��]`�j����7o�p1y�D�MG�e`�"GKmdf^���s������Xڱ�no�!V���GTw�h���r!�e=q.(��s�(���E�'&�w~����xl�8j��ó�WSSӆ!|�M�wt�~�����LLL(�����~Ѣ��N-HU3h���pp?�/"��T�;#J����@.�<ݯ�Fq	4�RRo��y+]u�c��|=�Eb���,���ڦ/-/-X�(<���T���c^����vL�9����� .�@�1arp� �1vƼn�e|�귺O��x�j�d頗ͽ��k��8�z��)�oV���ǼsNZZ�ѷ��~�ɣae��+�?�o���o`�����M �	d�U���3[[�Z����3���(e��ny{�ܞc;B$�XV1?0MN���PoJ���=:�Ou��)jX�x���xRr���S��mFV�6Rnab�7F�{�d$J�i���T�xo�zmr�B��Hs����1.�rVg���1H�ēv����,��C��=z��FGG�@x����\U!�y�0��q��Mr��	8��Z����^�EǼs��Pe�)��O(XH0�����#e�k"dt���_"�y��x `	/v�b��))�SM�tMm-���ٱh����u@� �C�Qy�� �ۏ�3�����8���71,y�����yh�ܗ��׆��xO???s�^��Ml}��h�d�]�H����l{2���^d�R�:�3��Hn驩V��Ư�4����"����-� �ج�kןx����Ex���o%>#��=�3\fȱ k��1�R{<��`��<�WYY�\���>�ݻI�V�.�-VKRT=�P+wssS�����x����Gx����X"�|����b�$��$���v}�������	Z����{0V�s��e��U	d��|�1��/J�a:&{o,��@�E$d��4!g��y��V ���y����۱�222�A�T���Ŭ8@A q���@�34��w=�I.�W��n9��q�<t=Tm�"�Κ"!z��S�����':�tXǭ!�޽���#+�KeJ��'�G�<G�XqA0/�́�Y�<G��H2����r갧�'��Ĥ����z��#����@<���� ����N�/C)f���" ��Jq�g��メ(�d������Vb�' �(��Ub���2�J���ۻwo!T��<��
��[���y1Ӳ�}xB�L�&�xoN	�|'P�+G�Ubq��C[����Qtӽ|�;*/^�ݩ� ����qȎ���}}E�b4&H!R�u
�=�s�'bLٝ��zm�!�� �O���qZj'j��䏲��O�I�T�{��3Ӽe��S衮���]:Ve��[j�
Y����@SR���	�"Y@ˮ�][�Ӿm�� �.�y�իWk%@z�&x�2)i�T�ә�۠�f���g$�tKU`�Ť���ֈjcЪ:}lх�#~J1u�����mPw-� �0�}�Mu
kT�R�Y�\h��E�u�@#V]<:�Yut;x�)��ι����X3��YOp#)����ў�/_&_HlC�V���[��Y��!�r�ܺz�ƍr^�Q�`��.��3����Ʀ���-CiJ1�2vLu�?I$Y�TQ�-?&�� !��@%y�(ݲ�p9�����}���PpΚ	����Z���\&{��kAJ��}ll,뻤�+D-N�<�w�ӓ���1��o�~v�ٓ	Z�[�x���	_�����`6`�4�r�a�<@𛾀�]x�]�.1����յ�T���Qǧ����ʹ�ndԣ�K#|ie���ӧӐ�<��nC�����Y����u
�لKI�@'?�����pI�"Us,��IU�/��0��o��4X��
��n1�D
�#V����0���|g�Ԙgn��Qf^�řr��>��Ǔ�L��ױZ	�f;� G�%D�p�q:�,Hluᐆ��333�����A�VY
�t����h��x^�L4���3����P�Ǩ�K��Zv�_*��NNq���x7s�!@��Y��%��:Յ���"��}��)\�	�h���a�uh�5���i��f��5;a�`ٵ�9�1�N��״��H$?���9矟B����^x@U݂���wɚ+������ӧI���:9�J(���
'W�Å�:����Әx�A�h��}��i�1�������~�����_�Y�.!v�Uf�}�V������d���� dO7��:͎~C4��h(_A�ӧl�;>|���j��!Ë�*���Y��7o��p6C��{&%@h��@��z]�K`CI��?��$%%m���6?5�lٙ?g��E��p�a��I�G����)ÞK�}���[./''GƎaSH,�p�O���8��Y��!��s�,J�{%�PQ�Wh2B��@��l �IOCB���c���dd��jBO��w�t��3�q�^�ڕ�Pub!��d]��А�(��������4�S�>�t,O�{.���̔�u��̂4�fU��Ie啃^L�}�T��8�F�T�� �n]up�.��Q�'X�����Ւa�d�r��|�BO�²1�">���`��Ƣ��q���O�*�^{��`Z@]����?��sƕ���"�����`B�}0KB8��2\S|��Ĕ��m��K �Q�E���J�}���*q�F��nEPT����Cpzh����;�R,ѽt�5��w-�,��i�#o�t��Z#Tn��� Y{k�â�L�|(�)j�xTΝ;���S��ꬥ�X��������&
�<+K�Ss!Ե�������a��pLB}�^Ksډ�Aĸs��*��U�4�?���5��m�ʴ;]���󈄄�^�����b�XO��7�=���>x{�	�F���[z'�jA�������9�>b�o�=��n�b�U
©�Gr�C�t3��pJ��p�( ������J
qm�/��Tz�Pqkkk$���&)�;�~��Fvd�����A-h��\^*�>�7�yeif��ƍ^'|��˘_�����H\\\ d��1.%$5�ne�n����3Š`@�?����c Z��.���2R �������0__�q�K{{{��O��EF"�=����{&��3�$-!T�;I���&�?|�(X������^��t|yߠx�e�Ͱ礝�� #a��djj*if��C�����S�ez�E�ҥ� �c9�d?���b<�:xZ�;?>��M�A{ɪE&��jj;:���/�̸4���ÞIzYjQ2�d����;��hW��L eY� �;_�����]K��!�wbN��ؘʈٳ`Y� �P�����*���;??��2��������}��˘�z@��V���/�t*.5����aO9 i.���5�رc����ې k/p�r�uk�����v�*#�k��W)�����k i�			=`}��Λ�w�a�߱�A}����*�"��i�u�3,*ߗZ����J��y��`���^# ��)�9hpS�J��pZ��|sf��\\�ӝ.�H)}�������EX}��t�UUUh��69�F����}��90n?s���da����#h�Q܎髒|���lO@���1�wGa���˗/� ��%pR2]}��!C��[��8Հ�l��"U����ðv�{]}��(t�h�	���]�^�����Ӄ
��4��R��r��nk�,�9@Ƞu�!��N|~Z�]�u����R<���ۄ�'���1V>!���}�L���w�����K�7�-�ɍ*��P��T�v�^���R���r҈����{�%4��E3̞���(��MɗexO���qr�oh\�ʓe�������`���i������u�[�QSu��>r�Mo��*�>bڒ�8pl(�v������C&P�"�٣$H��c���L Ä�{&A�����	��*�����R
��&���B@�h���]���Py�;��Q��Xc���%>,�]>|�U�x���_��"������
�� �B��~���&U{m����s���}||VD'C�^ e�G~~��&�u�%e[�Q����J�����Zu7���~������m!��z��#E+��B�6(���C�IR��V��[WAȡ�� k� H��22n�e�5��/_4��V�_bEkjj"��$Yi#$�n]��&)A4j�Zʲ�ZV����y�@ᮡ��/8A}����I�1�}� ���Zl%�X����FX�@�Nk�x����B�^�vP�8���M��F���e�.��)?�=gBK!y�K�W�ሶة#;s�l�>6��OȨol̔�z3	���4p�4�V�"&]$�}0{�~B�ID�'<2R�R�V�����FzK���f�C����p0��|E W'�U�C��#G�H�&�P�Y�_�����O������)��>F���?�#0�[� K�ד{�>ntt���Z]��]�F<8]��(z[ \$jaa1��"�% TP3���kkGB�ސN���/��)�]�
ɦ������@��*�:��6Te=�%�(��a�%�=V԰�U�n�F�.)���7lX����׾���GKX�.&hIS���k�*�������	��a��ӷ2?Nz�)�vC322D���1�����n��ǃ(ϣ}�������".����� ����H?��,����*g��G6�����/���p�����-3jt�h�c�1h���X���K���I?N���a/�*�ہ��3��sn���[ɾ"s?�G�鑳mvyc��`ڞ��Q�=�Wֽ���g�Pr�|:���kF�Ɋ�*�n��*���Bz����{�y�`�.--E�����K�H;�(~��K�+I�j�1�疙v i��*�>��e �c?~��[ �^�푔:t(���f���Y0Hc#/�7�>�+nz���QϞ͞p��VR����V�Q�7���x����q3����q��g���"!����
��JrpK]�XM�%PtK7Q�yí�L+���󰰔i0�;�S�IY���@�qǰ/ә�`����0��6��GY�LȦ�c9��
�a���~ժ�����;P�)�z�
+�)��P�~04�SmmV7�Y�]`��`bb2��[��U�r��iZB���k�����ڳ�@��=v�d��ͭK5V�q�|��Ғ!�V��
\]�2$���..�N է���a�&w�ܩ��@*�1�S�"�gH�� q?�k�`�m�N~C�͵Cy��3��Y�_A6��Oqh�<ZKHۛL�3<�x�����$����\&�9ϟ?�+((����I��T�cǎ��������<R��>QѦ���, -�U������\�3>�9�;�i�eC�v�8=��tD���@���NW�!T�ǕC�	��~P(�(�����������N�: '��6q��y��e ;!C���Ψkh��IK��c�� j����ɩ=Op��c�r%���ƾ��G�W�)�
�A��o߾ՂM?쀄��Uei�Kp������#G���H5�������Beb�!�Z^Z�C��}),,��GS���xlI5q`���.�N��N��?�8� ��`��H!;L�*Ctw�I5�%�(���k�	sgA��V)���6ʳldm��`.1 u��x����Ւ�{�2^M���^��3���LM�nD	 ���+�:5vw/��l�*���s��M�k`�<)�M)Q�6.0�}�6?�b�t�9����82�un|�Z�.'&�)�/�������p�y�LzL��ń��,h\��l�'�ړ�ݷ������ݻ��J��QQ㧰b����Y���4T��kiӭfQ���A_K7�-�vY�
o 0�b(oo�yOOO�sہ<��/�>��"#%u���^;BX9H�y��������Gt�N!�F�M��B��&G�,��`/\�_q�v���/\�p���< ||E~��1::�~L�`f�抃�ە|9o�����n�&P�� �B�WU��%�7"(�����O��6�?}�����v��H���J��Rrr�""##y}�D���~>,�d���}ڔ���q
R=]�O�`\˾��50ۍm��}P�D�W\]�Q��K/5X���V\_���
v��ʒ����j �j��
�x�!,�j Ԥa�Ȁ��uu��h�蕦ࠃx���-�S��5���L����[�#G���!=���+¯��� �
�bS%�i�;	Tj�ּQ���J#�0�q��pGggghB%
��ADMS��N��@�#��(ds��4���C�8����j|�����t�������MT^B3�q�f���+�p���orjۊ������)�v�q��C#��|��h�7o���1�E����2F����q�~zf�/Z��03E�;��&?�����o�7b�w�V�CM"�o�^�v[uR
���_�"�3�z��kkVF�R_]̱ofO�g��w�+��S ���ˮS�y���\��)O�p=3���r������R���		.�Cs3���n@��dKNɢ��\9�i�i�Q&��{�Ϧ�U_D'��AiB�2V��RٓgϞ=���A:�>���Xȃr8�W��:�'|&''��~���R{�y�@9Yx��y1�j����[,>%����~"+A�5+�n' �03;�� �����y���II��s��z{�x\m�rjQ|M���G�._�C�^�}���@P�*H:T�GO8=~��ϑ�LUrs[��,�+��}A�s�m�im7?7���e�^uu�-��-��ݓF��@g	�O���T�����젆� L^�~�G�Z�/�jԅ��GP����_��v�b��!Dۨ[fff�o�^-t����0�\я�C��5�N���n�����B�6�1���;�������Z7� -$�K�L+V��߾�$�8�ف�x9�okF3�A������g{�T^����n�́qJ1��ոl�b���D%�41II'�_�=B�"�;��*D���]Eq�ۖ�D�?�Q�T�_MS��;::V�w�R�0NOa]���h�ny�!a��K}��>6���J�t����%�ʩP�����p��*?�7p��˗/����!;�k�9�#G�a)q��J�}���1h����q��iG�-���E�Ղ6hμ��~��cqqq��]��S�琉
;�����eC������ ��>s�-q�v�=@�O$HF�����B�N'Y��䤝%޴�����d�psZ�KԴ)����s�|$�R�}����:�nq���@��W::�V]���PFVV��i< \e�T���� >���ۨ����S����꾀�----���Ǡ��v G��xRN�,/�,��?gΜ���q�7
�BM8i����-�;���XF���Cg0m ����_��qs���J�!w�\z���s�U$ �e����c��O���]3������I"Eq �f�����Eź�M??�� �}�*1����Pz��9!ʋ:\��,8�r����U�ג����Ԉo~200P���R��6��QI��W��MN��_>�<v��B��ɒ�/��hB�=>f�>�;��QB���ԏOL�K�
�T@�L�`}��H��vmmm&H] eu7�l=��TT��q�v*T���z�_�����$���zB5G��	at��m��1�I��ހW�^�+�M�Ӛ^:�/�ͤ6�a����ܶ�[+�D�+�|����g��ݻw�^�»|����ԓ������m:���C�Ӵ�F�:�R�TfFVʍ��/C}|@\|���!��YXx/������B:�weW���BeaYf=�5mp��f ������o B/�T2�wH:*���q�����}	2��+�䮢��/��$P׃x֖�ar=UFΜc-E�abb�yOb���o����4�X���W���Z*3��V@��[�Z���>F����J��|T�q�h�M�S�k>*E�^mhl�&��rs��K���
�]"���K����Q!|r�[Qz�D���|/�LW���<8�b��Eo�!�SM[��KK������>#E��8���Ń�Ν�iCx`�`v�!��!>�Бwi;�Whc�|�ܷ���޽;���]��(5uuG��'AW����T\O+(X�nll4�{Mރ���}�`����w0�`����zĨ���v��Չұ��]_����������w=ހ����&g�2��*CtF��r�]ži<�G��T��tR�z�t0�[y��Pa��7:TؼQ�t�%:�������uuuU���ZS���Bt��GoUH-;U�#��T12ꩆ����� ���lڈ��43R��+�?yrrr�6 � Ȫ_Y6l�ϥ	��4����ӓi �w�I� �\�{�k��,>=�=�1��m��K	G��
��
p���3�	%E�~;����A���)U��Ă����F��,�1!��
���軪�\�v���)j�oe���q��JG;;�f(�� ��z�>ԋ!P�S|�:`Y�s����IU�*-�3}�E�ݍ���S��i-by����ec�UrЮ�":
�s��Z��3G�� [W(>p8"v>|��ԑ#S�8lü9)�p���>��#��$iǨ�aj�I���5ƴ�5�z^}id�%���1��3P�	�?��W��Cuƻw�C�����T�ct���&.�������ԑ�4������"����:+u;���l^$ltuE�U(��z�����a���P ��;��H�ٯ�OTD�g�<����r�Ǘ�r~�������6%9����h����drS}�h� �;wޛS��ß?�"L�T�׾�O���4��G�؁C�CV����-��x4v���Pg�Ry��A����#�psS�A#SKhj�=ǖ���d�_�-�2u�t���Pe=1wȤ&=0 ix��&6vv�{�X�Ԧ��T�������˗� ̎ ����6���� }%�s:lP�|��O!�`moJ�{����@���J�'=�"^��ᬕ䎼�n"dJKP&7���H�J$y��P|�H�\-aQ��6��<���A��z�O����q�6��Bm��D:j�e�!}X�A�?�άm��ha���q-lhn�m��0���9T�����r�z�gX@���
�}���_`L��[L{گxD��pe��X|�&�q��v��b5��/�UPc�+!9��EJʈ�\ �#22?�,��
��pٝ���z�Z_tg�NH�ikk[p���RA�_\\܊����}��C��Ǡ�07���}"��Tg��Qd�Ӑ��LLHY@�l(P�Z�x�[������yiS^����h���:&!����Y�uӞ���Ԟ-�X�¥�2�ֺ�P��~�_y���kH�T��b�j9��F?	=��=����i;��]��x$+#����͉sA��wX�(�L���c�Ow������g!�(�|V���,��To���ӌʓ���:7n�*.�W���Ϲ̐����6�y�9�s$������H)B�J���-�[�ѮԀ�;ck;�W+7Ӯ�
'$h�ss/��*��� ����t��}~;���	��A�2Ys�̠C�{��(Zg���G'�@KH{=��Ϟ5K��.^�*�ƃ$��6�h*>!�A���<���/4��� �M�͝7�@lhhF �J��R1��6��J���n�,��(�2ɉ�	��̅���q�Sũ�*��!�\n*pE���>syyy���ʩ&�
��o뉘� �W͹���������[��m���~��� O"W�in�Uq�m3-Cð����)���Q8y���V�������������ZI�c�&iq�줤a^fn�I��M#�0����܉6�UIII+�Y�*TB�]�v���a_Z�lx��oL���UP�(F���`H#�� E*�8�k"dj#dfRPw�||jϞ9�x��5x����{�22\����qD+�X���)��/����[��f+�DBq7��+S+���#c��<s�r�(��3{1���ӓ$/�'�22��'��_�A	Jty	��&D�G�4���F
Y�!@̢�w��]{�Ķ6���Lqv��С����;�@��.Q�r3���� DB w���Yj!51��=�*7�ח���rPG�$�߿@^u�`����}^,����A�S��+3�(*���A�Nb�ܱ��f�����k{��(J�{*�*os޽��?�M�J�-y�\<�� v��v��m�\��
��g�����yPCT���-x�8W���J���Z�$�E������֗a��2��'ҟAm��ǩ��$���u=�G:ȸd5�G��"�*K6���-�z�W�NTK�B�i� ��>U����Dn<��J8(��RH�\�92<����(���&��Z����me�󅁔�$:J���{+� e��-"6��Ξ/))����2j�}[�ߒ����?E���J��1j�˞��.J�@�zfӧO�)�jFi-E�����o9�$�j��Q�]����i�/QR�?3�e\A�Vf��j�������`N[�0�z&}�m�����(�Wg|nџ�Z��:��H]�d�ޚ#��S����c�>j�3���/q{e����݈���MI�u�bbii�]��Bs;-z�;\Vz�&�g�L�����������[�Z����0������J���Nc�2�k��#T�ji ���$�]��	Ǒ��u�Th��|�Z@<v�X���磨�e��<������&%��$�M�+�T�8�x�а�Q3AK2��7��4qq��ׯ����n�U�AD���cJ\�5��(?�
���!_����z��U����eō7��]��������=1&�.����倔�8ˌ*P��kkkW��j�R]S#2�΃�k��m��i5*��%ǆ���]٢���M�'��2`�6�9��<��³����`ͯ��Qa*yձ*Yv�ӡ�� �Jm`E��Z�#����WI�����؟���t1q��$M�C�e||<�ҭ!5:��;A�!i��
�YT/��!��S���G&�?��1���l���~-�����<���n�fݨ w����Q����U�<����1�q�z{���}GN�
���U�u�P�0{P����B[=�6ll���(.��Aꈭh�[-�>5�WM&���� ��@=?E]��˲�����̋�_4B�^۔��&Q��TFG��	oI��5Xq��)_W0�	 S�@FB)�?[d��=������ъM��Ѱ�y���G�� e�WT���B9�ҥK�P��&&Q�P�ւyr�qk0S[W���)zzz
�FEy\��uM�5g�b��Ke��� S3�<n�Օ <��U^`}�+=�ߨԣw���q�Ň��Y����`3���j(C������������/�q��ߎs�A��R:�DR�䄢TG��$���ގ�hD�f��4��aG*%�������n��g������|���Ϻ׺ֵ�u?Se� z̲��}M
(^�'�|�
/�έO�����G�0:����Jv�m
���G� �8�C�ƈLU5��TyZ�9��oܿ:�I� ���[[[�n��?�/z��%���Q˂n+3=�����(VU�<,M:��������R����]��ON���%h�"$4]-9=}�/ee������B�F�9y�ض���Q�?���H�Y1�����5�+?��Ĥ��_��]�a��齷��}�(c�m�������ق;���(���T�BU$���� kgi�I*5L�{f��E��弄NA�WVΎ�ܖϨ�9��r��m�!U�T`Z����|�:g����T___���{��%j^5�*�E�f������?�뢱�_�����ϛ:��m��?<��O��o��y�m�c�D�_�w=rR,�HHi�����M���{��3��A-��%�c����G��0i
�u�ɽ�����}�|o;�F�s.�Q�|2T#Q�6"�.q��u/���hH�nlè�Ud	��N�	�s�.������K�-������l�k��~�A�m��[�Tv	�T����{�*��1/��������Cw���qɛ�A^si�D{�����ĺUw��(��'P_�zl�wvGX5 ��N�	�0욷�Ֆ��%��S��#�9�.���y�a��ԃ�r��u']���\��_��B.m���<P���i�xG�1%啂��T�Kn��=��n8�m/��Ү#o����%��ܮ��������F��,�s�o/+�>����/6�Nr�[�4�j��d��J��|"*s1[O!�	<�p��N|^c���|qJJ~3Pn�"���|{���W�>�	�� �IA���-��o�����7ӽ�dg�;��x�7ǳI6�ְ������G/t�ڬ���? ��ؠ��Mع��I�ؑ[[VS������5$�[��h��u%cn��=�+y���D�e��Ӆ�i�rB=a�8'�����DcC`g����?}n\�N�/�S���nw����S�����f
f�/d�]�Q���9a��8k~�5�����8�qiiY�����zztU�>���r2�x�T|cK�sA�܂Cu��Z��ʜ�.��:yeq1|��X�s�y�f�B,�*�/xTTTt݂4ؼqf�����aݖ�{C�T}� 1Ϫ�zt����2{ɠ�����>�e����Pp:u��0�1?;<l��!��6��L��.C]��'�7�k@�Z��z�M���vN»▄���ƃ'n�{c�K+���3��T^����Ymfk;l4���2IK:���Z�F���y���ύp�`�	�ps��ԥ%�]
s]��=��Y��Q�K�H���kii)�J����u��������e�e<�|cC҈����}d��ٳ�ڟ�N��7s�J*��J�JeZf����K������Ӧ�4�������KO�; Ȥ��8��+���[��OM����1d��[ތ�s�Z9zi��f��'N86H��av����{|�X>?'D�؇�g��z�P4��';�^�JL�w6d.?~K4@)a������/�`��,��	5��}�
�9�E�Y&���z"=DB�q�ev
���W�wŬ�y�Vf�M��o���;��4_��x��4#�6������j �3����7�p;�
�dM��V�=�����F���3;<��@���X�N��3����x�r.�	�"�j��WS7H������Z���>�[Z�L��=��~g���y�XDi:F��+U���l��纍��ɦRxT�M�#.c_��e:�S���AV]�P�V��]�r��~x�%EWD�qaa�e��>Q5�$�}�Z��<�?������8=$�����S�C��ts@+%�〖�&ݽ�"�KK��q�=�KA�����J�2�Z�ޑ�l��g^�n�mh���4�����q����Ǹn�&	C>��ի��Qi�k�IIIi�E3�*M����L+��5$���_�vU���k���zA���ck�|��h`U�0�m����fl�]�m߿;�C'˥����𷨩��b����#Lq5~�ܭ����2K!\�y͎1k�W_ÈY�~���V[KK���F�c�;cccG���_#V�Ha�n-	e��yכw�����zA,��b�:�V"ݖq�ۻDu����ļNK�Â��BJ�w�5�M���c��Y[sm5�ܾ����Y�[̯/�gX-*	=S��k5L�ŹС��5�ѩ�/����G:PU��eUB�f�^�5�R�M�"p�콋x"Č�s��f�8/XJ�[_��&Vc���	x�<bF��H��i\D��0�9p3���35�o\�κh�b	�h�>�x���Bh���b�22X|+�8��Bv�UO%�gM/��;|n�\��x�*1�[rFFK[[[�I)*I�y��*�����/0�M!=olq�|RaN��v(u02������ �N	z��>���엓�佦�������|��N�<�P������?}:�
�~nf2�����:��i�Hmt~��������k���o�ߠWh�qWO.}�hM��ː���h�p��ɞ�Q1㒢��ؚ',HҮSixZ��J 0Ay�`����W#�(ZM�t#Gj�4H�8Y�~�k�F����������F�'�8J�o%VJٴ5��#ص�X
��u�#6�ZJE��+>o|�}wu�hoM�p1����?�sƉ���W���7uu����3RR6�bb��|���F��H v>Gj�����
z6)m�~��ُ�	��Q�� ��I�f���y@�	?���0K�5X@�@aC�Axtc2N�y�{���Q����K ��B2��Nr�CCC�x�m�}z�;w���rw�P�(���#B�mm���W㫿@��~�Ğs�a?'7�vpp0����Q#<&���&b�i�S���_!�	���)o ����ߎ��G䈾c��,�I^5R�F����@�Z����)2K���՛�7��s���z�,� ���<��۪ �"7��W��0�Ar$��]��I^��{�C�s^�2ؚ�/���1��(��|�jg���}xn� B�Ϳ���]�B����Z|w|RxD�� ��Sa;z�^��8��E���|�Iȑ��/ �9��]��!� ��>�Yzy�z�\B�#��z�M�rvO��I]S��1+[�L���fϿđ-T$�����Y�� Ω���c#ȱ�c�{M����p
��:�����c�q�y��O�^�ih��MM w� F��E�&m"�n��o�MMM�ڶm[5�IMMM�W�\yB �����oNwJ�tP�rY%^��q�l�MN��^�b�;}��qr�]���y�8@�%�-�6�ܣG�1��h�c�4���ȳsTe=*y��� y/ Ȇ�S��NȒ�₧O�8�"��_�� 0��(�H�B����N#�וؤ�o���5��["�a�����zO�X�آx奄'�����uP��KֈO����N��{\��&���L4%p褰F\�r!We�ٗ-\\��&�@���V�?���?a���@�C�ù�7�%�)�
O����5׉���#O�43s��@���l<T�"�5������<Zz;26�]�0*�w�7��rԓ(�v�*+�탦	qY��.dGӱ��	uJ	'������� �!V����Ɣ����)6���c�(��m輰�)����zAWCpds����;�1ʤ��4�䎂�\�������p6��r|8�����oB�u�4�c��B�mY%�[p��98B�)ז�-����G�1>P�f�h"�ȧ��_-���bˈ?�p^��al49T8,�����#7-6ش�=vx/���e�m���䭚���vj���+�{!��˰����)�)Wa��\z({b�_�yv
�H��$]�l��i�0���Drd��F~��&�.�����̃f�ɕ��ϟ�5d�`�J�;��?��ڴ���
={z_tt4�����gyEk�����P{a0I���]
�fV�d*]B������V}C��c8� ����y ��<��e�_�v2���w��B����]뒒��A_O���´R����
��.��W�^� �zFQQ!G//�4f�.b^u�&]5�����>��n�>A�{�D3��7�Ƹ@�/A��du����u#|p箄zrS^OG�3�5eݾE�83 �f�	"�oA3 %���#�8z&p�4�5Cj��v�$�UUU[X�)��s㭶��K�kRF�
ڃhF�����5����=��ҕ��n1�v��0���PŲ(�И�����.�������'h�M}�c3(��|R6��@v�^��:9:x��L���`�
������ν��R���X�&9LL\Aa]��'Y�JāL���������
�|�T����T����P�[P0��hIE�Y�N��<G�ʠ��̸��QQ�A��ܾ�*�jhԥ`�F�� �`o�����N������%W��cIE8w$�q���� 4�����Q%m���kD[C����������&���?�:9�t��9]-V�S���O���эI%sk����)�{i��Wިg�kHf�A|���� o%�r��9H�8"��f(�nb��s|N��aTjyv4���b�I{7���ĩ]�=���Ψ|���Ƞ��B#4S!f[�����lH5.������^����0��ٞ��M����G]jG�ۓ	�a܊�X�!�|����ݲ����4���v������JI�������5p#|�_��y���Yǃ�W����Dk�@}{��}KK�1�J�y�N�#E����Qz�ƌ�{��馶��V�Em��=_� OC�NP�7���M ��KJNEEV7|P9X��G�N�#BY��p�c��!����T�;i���v�S�pW]]]���ӯSɧ_*գ��^GK	�tJ����K�.5'��sAy�;��K\��Hb��'���^�Fxꭋ�����A�˗a�(!�f�)ih����x�Ǿ��o�Aߚ���@��G.=+쯡0���ЉM7Y>���Q��o��Aà���3��#��W��[��	'�jio7t��K$�"#���B�蠭*�A��y�tP�
ı�pC����@��<����6��@���ḥ��Ī'{w+�7"�_��O�"��A�l��^@��KӴR�j+|�"����s	��H�������w�`�ñ���'O�	��d�:��2���dQ��_�P ��J��E����QQA����Q��_i;�;�������8���0�p�22b'��*~�Fm�7�����O!ި�C��r��`���OI��
�]X�ϖ�\�?���������
O��Q��1��Gy��-|s���|�'ළ�}�?��d���Nk��4u�Ij�"�j�˪��n%Y�D�.=�]��;��������,�߅\�b��RUQ�v�À ��,�έ�*Z��J��]��c4�s��~wwi���1�܍��/�-��O��Tg�����r�f�M*U�ژX��#[�U��Wtm Y"��ȑV�1G���:��p5KԼ�}�v�g����c�z��o���O��wUB�x���=��qqqe�9z���F˱�R��Ցk��][���a�6( ��Z�Ƌ���E�a����dq�΢��Q8�ic
������p3%�`C�cN���&����y	��[�C�f��Y#B��,���+��xW�����������/q;�>:r�%υ$�-�p���hڪ�.�)���|�U�~�t�˨�ïtD�۾���s��D/����m&^*r������W�ᠳ3���,Fà3S�c�]�Q�6�K�OÚ�zU��r��"|��^N�N��J��Z��v�'GO��`�V�RC�<�|�͠��[�F��³�,HO��'�QqD���S�Rô�N��5WA�:��@�섟�c$�F�������>~k����^̐��-�G+4�_��{�I�^VV��dXGR�*��3�'���W�[�E��0K=���o������u��"�#<�P����%�$���9j���8�\�)�9@���/�p?�l���:|��2���zmz{��d��8��!�k�,+!�d�x����h�@���ts��Ç�e?�5��.JHI�N]'��]ҧ3�
��U|)��Zr%̛�ؠx�r���y�Op�g
v����-װ�j�R�E��z;;;��x�C��4��>���<>*k,�wVhn����ts�������:�#��~&;�k܊��+l��ۖ=5E����%�8d���z��o(�(#�af�O��\�#�W&n`0�˂H��'C���9�,u���Ӗ��K�76�[��nl�&̍o�!ͪ���D<�=@9%���X�c��Y�_���O
�d�{���1��%c�Nt�����s���3��]Z�0%�	�[k���ց݆BW�z
>K�/ �t;#8����g0�/��`\Hو�Ʉ���\H�d��:9�GguÓ{z{�е*8��,-�G����*�w9xm[�UZL�d�0M���XW����k/�}|�9v���wEk�줋�ǆ�[X�����M8D�~�h2f������,/..��/��Cl��XX��*u�5�u�[�������3�!D$�{�"��Ý�h8%�ړ��r��s��
k��a	�!>����5��]v��_���(SN��.H�=$����?-
,��0ӭ]����S��ٵG����h�*�8��u����"��r65%���n���U,lޘе�ʝ|ŎP�&1��V,���)�G���E��k�ЉOn��|��^<(%E%5�@�9�l ���6��bI$} V5�Y��qgF�������0d"&�n`�s��Y�x"�p�s�b��;����E���K���b>o *��W`㊮ ������%�'�z�9�O�[�����v�ݼ�vd�Xb!�ۋ)Oe�'��v׸���	�Q�>��d�iral���V�������ct��g�ȋ�}�PGl�E��MI�9��'��o*ң��x+vv{,Xʐ�a��g������X5���^,�>yD漂	� ��t��b�x�Y�5n����v��&af�E�����y��m~� ]-�ޅ����<��w�L7�Sh�3�����ĆX,P���J�T��R,w;�Oc�'���ɠ��q_� ~vn=H׫�I��酦�;4�p���R(�ER؜: ��֍��&ڟ���bF�Яu�t6�Fy� ��>�����
�VDB$��b�����B��d�+'n�P~����Ǣ�֔c��K뱛���Ő�-	�'e8$ T�����"3I�<������s+��m�ӳѺ��a��`3�TZ�F�B�R�,|'((��y�/�
� KG�����Q��!��t�7YF&t3
>����
��TCfCB��K���)����3)���Z��v�H,O�A&ka��czB:e>��c�~Ze`Z�nߧk2�Q���V��{��ʎ_�;~���-Jm�+e��%��_�hZy�aw��/L'�f��m��][�s<~c�"�A������c��Z��^�y���Z��]�v�`����2�d�F:(JKǪ+�U�-���k&cnL�sn4~^*2�<�B2wN�(Ȯ({z'��[˄�Ol���E�uY�*��ܷ��`��; �^aw�('�*2�6(J��P�{j��=Y��׶K�T	��\̨�yP��"���0�	,L�0��A6���P�n���%�k���J�'����u��p����k`�ƛ�z֭��T,���C9�� a�-��jXX�ɡu��������9?��#g������C[�������'E&�N�����|:��zn���'�`y���1.�i_1�P���G铴�ie�{����ͱ�@;x�"��`�!Nl�9�}8��~�F5N����`(_���-��Q*�n�*~��Pd��n�I�4�j���N��N4�\��u}��[`z�'�˺м��ƚ�i�SLr1�r�=e^,��8�;�*�e��M^O�x��˓���L&���e)��s�����Ċ�z����>�#���nxF����qUBk�-��[wͼ���B�݃�i�2q�W�����B�a����(�ޫ��.��w {<�󯀖9j�~��C47�㡧�CK�65@�ͣX��`wHu����n�;&2XC���߅���JDkx*LW��^��Y2�����  �b"|`��M|���V� I����m!�w�ܙж�~kN]�R���B1�ə�aW��ħ��!{*��������n�����q�"ڶd��`��7�����0P�&L��2=w�䚌`�ͬ]w}}}9�t��B��z[�Ggx�����rH���챪�[L%]��~��c�\B�a��ݤ��g�}�HUi�/_ᛛ����!pMd��&v�BvP���� Õe#�X���G��qn/���#��� �����W�9;�̽��f�S�A�&O�3�˄��DH#C��i6��򹒯�)9�Z0��K��ȒB��V+��\j�ݸu�Փ�?O��=��%h�Q'C���E�̍Aڂ�n�,C�R���-��{��Xab��v�<�/�{���#O�6�-.�D[oW��=;6:q|,�6ۛnT<��L �J���={���ңpIC7<��~ya�F��Зb'PM��g�+�U/x��﹦�(�A�aѹ�,#�p1{��R�xZ����ʮ���`pa7N&��?Lv�|�> X P�]�ש�e�l�Z�}_a��� ��!�\��\Ú�3F��.��F�v]�ip�u�!�����t��nd������q��R�S!H���3���{�����8��&�l�\qx���r)�q��DF�چ��A珮���û�K��O�;�o!ţ��$oʨ�$>���7�YR�}����
ѷ��� ٥=]B%8r ���I�,��2��رKHz!��oR��}��@>|L7�/��=��%�J���>�{��ڱ�島�.޻�
�U1q˨����6]����9U�8y����qcK�0�bǈ�,�co�{����xC(L�P`&�#�Τ���v7�y��WQ�o��/WM��jl͝gEK�N���v���pQ^m��'�K�YnȜ܎��S?�+��?�s�E/pi�$ab���Z�7�ї�<u(C&J��[s�rKmv��&�1����,�aDb��'����9g�zۮ�VI)����~�?v2��ӺR��A�V�0��Rz^�nfk��J�$~E��/d�ކ_;���,Zs�k�l�<ޮ<�V `�B�kW���l�&k��Q71���{��u�jۈL}Ux�Wr���X����T2mJ���4T�Ԕ/���z��B��U�3/g/�kV���`<�g�� {��Sj1�Q��%罔Ґ!scX�W+����<���F4�R��RR�����{~{��|�~~���>��є��E�!��C�j�x퐏/ݤ�������Lf��L���m���X���Y2��E;;�o�ꬃ"��ܾ7V��ڟ��م�4�D�ѐ}���S*	dF�P�q ,��$��ŋ3���c��Y5�-R=�Xl�����V�o]���+�l�]�B�5<�e�Q4�
�f��[	KX.�/
���eI�B���(���P�'�"+��.B" T�bz��^rE�e`��=CDU�h�0ǃ�F���aU�*c��At�7�ևi�b�-!U�w��Xg�i_xd��T����{���,�/H�Q�ɠ[�Փ�z��Y�E��a"p���W�An������?���c�E-�.6�B>��I�pE��VV��@�=8�P���)� ��kY�
�@�rz9֛���B�$�Uf'K���T	��"J�ޥ����}�O!�� ;�b8�
�*�m�A��M�#!��Ȳu���T��+;��e�@������_ L��µ�Bڦu�T�R����s�� /�r͡�N��6Q='�u~XQ�����
+�&�j�B�4�?��Ȁ	1"�(9�PA�T�!��ν��4ϱ/�h�:��ѹ?��c�o�����E{!������-v��Li��MW��rB�0��u�>(���.h{#]�K�+����;�wuD`����E}2sEk� �,��ߚ�گg�"� 3����]&X�T��G�#3�N�Q&�E&úU��@�����E@g���#�Q�/���N�)�����K�ݯ6zd���8��uT�(2l�ձ�ETok��(Ah��x8����Tg�|Bi�@�܃���RRj%�F��l
�LI����-*�����S����׼hR2:�p����\B��
})�-Q5�	-v{������D�jb1�x��@�j�U�$ZD�kAFYꉄ?}������i�R�m�SG
$���_�m�F�L��2f㱵�k�s?o9��M�"O����,DkM�կ͞��P����&�*cn._���<G��\��c�<�E�<!�I�nIMM��D0�<���Q�h�/7g/���Y�+̣��A8�������� ��0(�z0h��%��s���;��ɒaø�{l�C���=N#:���d���'��̴Q`�Ɣ�@LI˜�Vf<Y�-I}�S+A�Vgy�'��*8rc�Ҹ��}(�^�-ND^pشdk���Κo�?X��{e�]�v��]��s�[��7 ��s�a:��Km�3��D��M��g��G���eB>�a��n��<4�;�4û'����N�Ů0�#��b$�R��c:��zU}���6����]&��{�����Q�g�*�G��t.ݒ�_@�Cz9�TjFR(`��y��@�Co� ��y�q[r�0W�٤��E(� ��Bor-O��@OG`p?\*�͗��t��ڄ�����^K0�-~u~�&@b݃����H����0m#ݥ# ��Ijcd���vy��Nl�XS�~ '�vF:
��Nё)�
M":�u�[7�x{#��ח��d{(5"�;j�uCk��j�A,F5�DÖ!8�uk/���]y�))�"����XE��))S.�IX(��'S�ڸs���9���8��$��b.p_���71�o�ޢ]%ɔ�/g9�q㑰���t��F�}݈��j��	{7����<�=��6�vԙ�a/�W4��9�,p6;F��,�NY�L��C�H"�10�gv��Ú�yO49��8���W ��A�1A(( NOBuP�����1����?��1�v#Je�<��GO�B��i :����sB'�2|⍫����GE{)	���$�8�}(p��%�#Sc�
(r�ؽ�#w�E���4Me��
�Η�A�2����mB��!l�aaЂ ���,���3�9<��:��C_�f���`7�\2�RRp��O���޽Ϟ�>�Mݣ4��� "\O�B�9pO�k���^3��.B���M��$=�u,��hc��I���K�J]J��:� �މ�Ԏ�[�J�ch�H:lV������}[ی�v���A���0�ފ�X�� SJ�	�_�2SR
xM�A©�f�	�j��=�Qs�4��E�0~g�&��՜�;9g�L��EŚa��;�Y2cA� vږ���k���,��:c-�*T��^,�0�"���ee�+6G��s�5'�k,�x6�f-R�&/x����~�s�>� 5q�����@��X��Kg�B�U2�5r��۳̀�t ������ބ6�̧���@v�9��-4^,h�����Z�E���uFL�Jh�C�7%C�L �P�!��f��6D�B�@���|�w��*u��olđw��uM���9��"Jr���[s@��A��f�u�ģ햋X����7/L��#��t���PJ#-������Pv#���h��b�M.�T���If����9΀�KU"��<R�5�2_����W���P���U��$���e��A�i���~�ͬ���	�̿At�g�vE��sT7��0�J2�g@���}6B�P{{�:%����х� ���Ċg[�%��(̾�rU�"op%+��-Q��n��* ��틸R��1!�ъe���u�5�]�$daiQJ�T9o�嶍#7��3fDjf.�����P��)��x�&G˪�����	UHf��[�ѭ�X*/��)��U�"/
�1��t�zz
j����<1)��lX��"�}_���}8Fz�h�S{>Ta�����fe}�@�O#Q[��ezή5ǜ�n�[�B]�P�2��|��xb�r����/�M�TP���Ix�m>�����j��<�-�2К*�"��J�וރBp��9'û���U�����s֯S���'>vY.�S��U-�K�F�����Pl֧6^�~Nv&��@���*� �G%��{y�>A+���i DT�F�����Ŋ�s�Bch��.6E�1�l��{�ӧH����&��:��B�e��9T��í�|�ڨ�0�$i��:l�k�Y�o#J����Ek�����b�B��:����_�]h�X�y����@�g�Ȃ���ݪHSl���r�e B��nrx�4�-�3H�B��]��HI��慺6/��+e��łJ����2�f"��@�+�T�����N�-����v���O �:��-��}�j�3�������AJ���	�h��$^O�h!)��>#� y��+�Q=�ѧ"(q=�[��k2{��	�Їӭ[��n�ГAbx�	b8 �d_,9>8\s��ğ+�px8<]�^p�93�!�W`>P�򂦎Z���\�(�l׿ї�T#voDy>s A�Q���,�t����h�a��&P�E99�|6
Xb�����XI���ahF����@� �5��.u�FyU�$��jbà�7�$.�{Np|��LFX�ٶ�|�B��V��A�G����wxRJ�X���GM"�����r�r�?6�bM��tI")\��޽��ӈ�h1��R�T Ha��ޘ3�͍t�DK��ܱŔ���R��H�G��[2��<����yM��m�6�[z�B�߀-���#���W�h^�o&��}Ȏ,������q;.f��q�� ��RR����޸�R��PIU�Rk�YpǸ*��.�����7f�1c�h�}����	1P�11_QfWd�Z	P\����m���N���q��Ե�ի���ߖ1ӝ�擲�D�KG	��@J�[(�<�J�Ғ#�8��/�Z�f�@g*�j���`��S�iG�q���z�������s��j_1��:�CS%���ja���T|u<8\@ɼ�a�y?��M�%DG��L�_������N��Z"�&_��'L~��F�H|ˢ2�xwi[�W��p�_(���aY���w��Q&��ZT'�{[������Q(j���k�������L'�b�h�ƴ�4�ˍc�4[Z��#ɘ�����4�m�S�2G{��%��d�����"Cs��ڇ#8}z���LeJ�^�'iR	<�`xz��ׇ��mff|9T	s��k��D�7�f����ʶd�4<}�H��baK��\ZJ߈vK�.D�<.�Tnh ���3+�{v*E�%"�f箯��r��U�!(~�����":�()����9;�>Fr?߼0�8n��+��{�Q������� �[K$�ؐ�oAD��]�F�	�횃Tx��X`|�6R��'����4��bv��4 ��O����z~j�ō�A�U7̝D���ǿ�datLdr�G��k����)@0\#9���$z���ȉ����KԀ�/P)4� �K�K�d�����w�y������*ꤦ|�D3KJIф\SD7���-���I�d[O�PAUu�Fy΃-,$���1t�[�r���XE���Đ3�m+)�ǐ�\�C�^����@%��d���(�aX8��Y���yDKa�y1�⿹B�&�b��W����A���G!�� Q��B��L�Њ��#g�=�u���ۈ�3K(cÏa�d�g��$�	�;*�\F�LV�:0rj�O/O��Ff�w���&��U1/H.��qr���Nl뱡{��q�oJ��i(�@�J�|⍠����O41��v�f��e <�P�n�I��pBV�D�#j
Zxb�W��@U�B)J�fba0�XJJ�o'^�DB@��P@�̡���������?��ڼ�ī�H��}iD--BH�kt�5�x�K6�T�n8��r��F��F��3�-J�) `���ū���c�"M�j�Ry0�8hi)"pE@��!{k���/C�ՠH z�ӆ��Ow��5�g��l��Ql���1�)y4o�_`��|�B)���;�Ġ��Ea%~���0Ū\�:=E|'�'��P־|>h0<b�t!n��<��n��%��k�~�
۩m��aK�����ܡ��	"��������b�w����k �O��JZ=���-�Q�3,x����\fU��R��%�]�-��ù|�Ы�gx��e]G��aySD
�Z�>�yM���P����}�d�úsPH*"��&O��z�l͓���+Nq�{�\1��)'��_L��=�ɞ}�����V��Ő퟿"���T�SY� R��Bp�a�}��	��AaXR�Z��y{���"���c�D9`��N������tþg�#f��o��RgO-�1�NhLkN���6r> N��qWP�����X��b�����XX�^[�Q:�B:bhI�҄�t�(��#��w�?@\M�nr7���>v�!T�A>�.�k��m�4{^,�c�� �?�AJ	�����BZ ��dJ��&p�W����R�c���6�2?�H �H�)
��
���jQ��XzF����M���V��c�T	��(�P��S1/��+���V�S,�(A�{*�p���Dk�EQ�?B�C�,D��GLiV��^�i��A6�ҡ<A9er�J;1��j#��E�Ƃ�.���!�颦2���3�[|�d��=5��{�Q>�����n[S�^��tA��^�!,f7J�����K�W݀N���X`���Zrü<6[c(h����Dx��(X��%J���&��f�5�l5'rf]����it�i���!��1=T��]ʓ��QL��.���rSj��]�Ҏ�Rw��J�Ȃt���s�ʮU��s^�J�ɡ�����k�x�)�J|��Mtf;��b�E�ޙG9|a��Hp9��̮4=%r^�5g^M�K�$L�	���ל[�����\��%:� -.��%z
������e#d��E�����܌r�5-:@�7�Μ�G�&~�76��R�0�Yy`�M]����\)WVn�]�<��_t�~}�.�j���̶�α����U6I\t�ٰ�@4�/2�Kп�Rb�Z�7F�7lw�8k�3����z�����~�9_;����,�w^ ��m._��I�P"p(���3v}����{��p1{Hمr�RB�7a�'U�y�乙d1�g����M�ްz�w����hhTR�2Q�=��w�J�M���1=;���Gل��T�R�JN,�h9����I���va�6�'�#�؄�~��k2��ƶi+�	a��J�h�f��Ϝy'���5�XC�X���2�f}?�N�k�F�ܓ�_I��N����u$(���ޙ���m�w?i���1�I�Y�
�R�[C��0��ӓ-����~q�����fʦ�Q�����,�;*�/�h�{>�����a��KB�oUa��9���:�O��f�3�_<Du�������ϸ��|�U�k��$�;%�z�~
�)ﲦ�m�f�="/$�\;�y��>x[��5i��b�x#�҈mG�{�'� Q��}Q��DW0}�~NiQ[����oJ�s�)�?ij�A<���%��B����.Vi%��Rz�Vq+nr�9�s2ւ���M�
?�0� ��<je݌�$���0S��ɏ�D�����<B��-Mw~���O��]�J�_�F~�_��[���[��[�i.\�W��w��m�.XDQ�q�[y�H�j2 ̛����Ckm���X�b�:��I}iz���Cfˤe;A��or�c�f��[]uߵ�L��g��V�~�]�f��=>J�̇���W�g��j![,��%a��o�����뉕t���Vr)=���1�1<ہ���V�AF�;W�u�'ӹ�@��:p�*��4��;���ۤ�9�T��,����g�Q�{h�!��ε�;L��6r�
N>Q�~"x�r+����H"JYb�Ȥ��"�������hh�ۄ���-Ӭ.^X��7I�d}߲L8��8���������)p�9>=[��.d��UEe2/��������?S��f�m��0�zb�t�~�����؅^��Hp[�9�����\���T٭D�IѾ�%��ғH�4U��]��E�$��$�$�r��땢ͳi�<�\&˰%���V�%��.�;�%��z�D�(͸ub�7��J��O��ʡ�>
�����z��n"���F�OYm���qZ�Ή5�-�άƄ�X�k#��ȘQ��5\"D~��:�}�XJv�d4c2�&�ˈ���W�d�*¸?C�������7����`Qݜ�$�;�Efx�6,ʝ�$�o��b	�#���]Xk����S�"?c#d�~����E��lլM�p�O�ƣwF'l�tRQO���B���½�w�p�!�u�c�O1�a�CG����Y�ad-`��գ��DV��"���D8*�(5��5����b`�f_�[x�N譄ӎ@ �W���/kV�m's�f�b�0�9&�-������#)�S25��I����\�.U|jIg�����s(S�����\�b�P�	��i8�z�^��T���{��2�M��\\/�0��h�Á^�e�w~��r��4[j��=�8�Heb�ף3�	�G�,�Z����6�,)H�N*��3����?[+�"R<^I��d �(����*�����:��b#`8��⩋B��a�p��)��h�Pb(���D ��؀�Cirb�Q��g�=�2D=rt��k���#���h�Ϣ(����a���ZVc^�lO��Y^@�D\_�����?��̦d����2,V}`^������tl��JG_},8������l�p�A�Z����Tw���I��`˻�)���֬N8��5�L|�k` ������#�qwҲ���2LC��ېc��X�	�C���74���^��<A�Epwܖ��� -��J�5g7,^��I_Dq�X,���'��*�S�>(YX#�!��˧���'�7T`@���ԍ1���!�K��*ޤ9Pg7k9��I�h"O��  >Xߪ�d��ѝ�E{��t�oM���=����͘'5����	�*P�:ݠ*�Ҿ+Ӿ������у>���42����X6#[r�=��܉��zS���/醢�PP���砲�i=m�T ���^��y���f�_(�}�I���
�ӫC&���_�1G���w�7D���Q( 2�^��� 'Ǒ��"��-b�M_b-��'>0��h{��e���&��w��#�n�6�<Z������UNa�t�ee��}Q�T}�̽����/w[�gK�R:�R:��6�q����D�����]�8d.�Ec��R�葄C���μ�
IN/�`�9<��`Mw��w��"����M�*'�
��8�m��?�l�#��Y�N����	isB��4�g?s�vH�)� ���Mɇ��w.�����s�H��-I���PZ���q�<�N��K�͠}@o��v��)�"�KϪ$� ��[HeS��b弦����=s�7
��Џ��ӲeC����>y����2��TQt�Џ����x�DVq�V���&������1mM�yх�7uIs�^pb�6%�.�w��b�_���5��ˇ���ks�c��0<�`�������zJ�K�P_���ғV֣ϖ
ΜE�_���#1�]��V��hY�װrm����������d�;i�*�̠ٜ�Z���FSk�o�Y�,�E��i�P�saY�3)��#�5�#^����p�]v�G�x��@X�+z,�E�b8ڽ����k�U�u��L=>�����M�@|�S1{�'��K�>�PZc�_o�����0�w=�����#*}g�� !z�[����m�洠�E� �C���"�i��C)�м[m��כ�V��E�
�)��a�䂇�	1��?δ31o��cV�W��t��>7=�˩Aˉ�Ik,�I��{�I=L6���	q4@[:�>��&�ݦ$w�#S\u`���L^���^`VG���i�E�{=���ށgk�(��n��_9R�Y|ta�K3b�(��2-Z��\����#V��"�����2����RP�d�	�ю��b�W��:7�cRЌ�AF��V�[�C:�?��@W�#�U��s<�'���_vOJa�W�z�����R-�w;U�|�R����
����+�2���	��
�t�c.?&R���*"e�u����E=G�(ׅ���Y�����P͎�&�T'9w��awH"9�����J�ag���1)��`=��b���`��Mj���j�䏢7�c�{TF�t�ؕ*���+81!ăH4�|�%S/��������g���`�M�c1t����=1�Z]�J�m�E��ߤW��`�0>t�&T�d��Af�&Ν���]��a���q=��7Zf�d�AN�t���B�o�:��?�X�D%�%��:����S���g�,�X����#w'�Vj�1-IL$��6A��������� j�&ws��9���W�3f[���T�:��0Q~)@~�͡o�Q�>�E>��|�7��yơ��(�؞k\?q�G��
4n+�B��`�u�"~k��2��=�f�����?~:W�׏�Q�h���%�a08�����.�W�ὶ��7k��>+�t�����X��}��O%��2�r�I7~�N�O����n� ;}��l�S���k����s%��9zT�2�<m?��!)�u�������wI뮂��ڴ1m���}R��г�-F�"^S咨�Q �X�� 
�(@�-�����Ǣ��f�i��齄�d[1��庣ia{�FX�����=k$�pjf����A�a$�0|��""�B (Ķ����Q��,�Pb�?2��)���-���tP�^��&��<8���]��A��5Uts���tG�L��v{"4��{».�����׿�`Q��U0ڿ��-��}·5ҷ�J�Yq%,��`�G��cR�7�8�L�u�b��=<w��?������y7�}��Ӳ�,,���Do\jf�fj������L���7(�u�!��.l�ݚq��2��XƳ�d�8�{v�H\3��O��n�%�9�%\	�ɪ+�L�C����m&������E@��*uT�FS���p�2�x�)��$aV��]2OZ�k��Do��e^�#� ���=�a�0�x�=l�JZ��т7z|�C�sCF���L�/Y(ȫ��wܜ�]\�����/��K�"�m} ���4����?��ݒ�iYJZv[/uX�4��q�d���)�C��W֗m'��!�60f���y���,�9�u�x���P"썰L�s<v�-~���W]�{�Qt\��{� ��W��}+���6��Yf�%oN��C�8�	�id}ѩ�|��Mq����~��R�� _���1�O��"� F�lP>��P�K���UH����4�{V\�%�2�/[;凵��_Hާ�}���W�^<�G�����iO\3�:�i֓*_�hį*�y!gxs�2��iECa�GC��8�������y��Ө����~���S�%F����ע�zCsZ��l�[.J��K
���7�e�.A9X>`��1߃=$_�(/_�jݐ�鈱��2��.J��_�����x�����{S7ѽ����ݨ&K��n]*��U#�ܡT�d}ZdK�Ie)B2b�F���${��[��{�3K�������}�ky����9����u��R1�Y�ʪ�.��$:���}f"�,TƗ۬��#�9-?X�ً�o���S�ş���q&���t���P�{W>]x�25�����Oz��AYP(:N���h/x�$z` ���q�� <��??��� ��h�|Q�XV�I%���)?�(V��	�_��\�ĬF��g���aF&9�|n�������0n�~L8n�(�sUvu���P d����4�B�8MQ���v�v\�ol���[�;��D=�s�`���\܏Tt@����}	��,�|g���2F��q!�����'>L���v����TV�3�ƶCd��C����?�3D��%k�Ь�2-��;Pg��u��H�1�Ч��eʔ�U�언�1�m2,���pzɇµq������:�8������߼�i�A�[�"��Ҫ�f�	S�f�q$�+��xm���g*�z��v{o��n��|�_^=��;%,��(�J�A-��7,����)Ѵ���V�zAƈ�����X�U4���a�{�[���ŝ�l���h�%HA'Lx��M���p��%#���8ytY v�ջ����_�C'���c;�<h����vo��,���ogw�J�ݵ�s9�aK�%�����:>=�:���-�����Pʏ>qU�;���v�H�7�����r�[T+�e����0
����.�w��\�P���{]h {�wj�R�+b���8��^?xP/�������\�	�Z��oމG@H�N>g�yn+?e�6���IGcQ������ߏ~��b�8ˇx��(a�2�쁫x��n/�����~�7���g��������;�xIc&�(�j��5�عk�Լ[�e"l��3J-2�L��1�TlDT���@���&s�k�;�jZ�'�ۖo�#�$��#�AU���-��fN�tɔ�Gզz'!Q�����|��E�<2���]F�O�nq�4G�z,?����Q�)��C�;+2�=�]�����_4On#|¶rHn�s��<�S	��Tns��<��/�����e*�S*얃StK0o՚��M�y����v'�a�:��:Z��j�Ӈ2߾v^��2�1�4��?;�>�8�B+ϟ{F��	>�6�dՄ�����0!��~�[�H���6k[T���>Rg����?���fi�� ��a�Y�s;�~s{��Դ���/読���I+�������\W>R��.��6җ6�o�����t���hU-�����'ET֨�%^js��{3[�]�r����G!L�$�J7���fq����
o��������2�[Y�r��5|��~���'ܡk�@g/�Q�^��)�K�!�v��mxT��d#F/��a>�������ˠ{�!� l�r�@�IEFF"���K��/>�\�?�Af{�31
V�UQڣ�y���x�8�[
��q ���?����n�H��Y͟ϧ%0逾���1��X��8�!��rC*	~K�_�t��
�'�����\��g�&A[�@�ۇ>���`�F����]��k��`����֋h����!U/&8m�^�88Nw�p�=g)��EĞ䎛��1��{ǟ�=Ϩ��Ƕi ͡=���v�-�9�Y� _�:iL�Αr������f�8[Qt�G�
BԢG(�ooq�(�4�T��w���ř�JrV��页N��{��z%�6_cCuh� v��N�h�5������� ~T9(���ufF@0/*����F
�t��Cg��u/��Ƅ^�i+��]��̞�����w5g�����q{���n �_V�`���}���/{�C���K��j~'~�P�^�`p�	����}�J��x��hi1A���3~M��5�?j��8A�Q:������О#����3ɝw���*����e4�{����|YK�xf���ȂA�}��5Z�1�x�V�{�x�ۇv��E67�-�%����:[3���
j�_#37˖��e�A�^љc��+|���绅�7v%�Y)�H�]$��V\Y��;���"Έ�g��s�����.ϖ��*�f��:W�3tz�a3V�b��
[}'�7��~5��S��+��w�Q�z��L�Õ�:H��i���?���v||��l��v����3�W_�z&����+�܋����P�D(��Y6��1`O6�w݀�1rɺ�Z��33�=�M���WN� �Aɯ�w��{�r�$�n;�d�J �����\�Aܿ��n�7JH��jqlɯ��ۆ� x�qr�3�����4��,����Ƀ�3D�V�]626>~�g�n�oӳ����W0m��6��ݼvp���qr��[��ttt�<�Q(���5�y����8����3բ\KG�[�7�����{K�y?K^4�w�.J�r��vWa�%^�٭g�Nsw�q+����0�?{�`y���Q��MSS37�_��VC�d��Y6ZXZ^ o :v�hR��rf���������`�#��K��p]H�Dg
�:	0�g�~@O�o߮����F�p|LR�q++�����y�h)4�/���7�󍊈�TV�I��T)K���mE��K\Nh�G�`544��/	|�?F˟\�����<�
cŅ��w��޷�m��8,�:�TW���a�`�B�~󒕕7o���<�������^^l�nS�C^���o۶@E��}���	��U#��y�ɷo��z�*�T��ed��)����SYw!�A*���@*8�^8/wYp���}}g�A�&�']�2�!L�"��1�C���ʏG�C�y�ոp 8��}x��?�g�� �RR�{)z&jaGɖ� �l��߄��%��,�)��I��W��&�xOu��9X)ӌ?�zwo�9����oPZ�=�o����
W�kRbl8�~t�¨�1�>������k��;�	B�"��ޒuGS6_�)J��g�4F���8!2**%��7��0j��#4,l�^-�/χ�� %F���W�<Gg�j &�2(^�_��R-7DY�~�����ᖰ.���h<D;��U!l�0���q"��~��\��8��Q¨
��c���22^ەm�������c�-j�aP��nn��E-���p$�0�wPY%nL'�	��vZAf=��+%�}�OM���7��-��;x��Q����e~o���B�@XVm5�H��ZX 儷�zSB��x�!*�Ke �Ƿ)(�E�v��M�ܯЪRüL���r����8�{/hT�h9��'<�PSS�0� �Z����7�4l o����%^�G/Wb��74A:��^�y+-%u֎�S��;f�?��+GF��	����N�M�aPP��nѳ�C�po��R}�֘�ty�ѝ�B�ah�L����5R*~9�V}J��hSj?��kU��P�}aM� �DT{5mS�Ȧ_��+E$Mm��!Jlt��N�H!|�������w�⇄��)�� F�'�OP��i~���+G:::�jy���NKo���ĖE�f��`�_�V�+l�w�@��w?_o�GRP@����`�E�{�:�15~H���K��|��xzf#����'��֏�w�F�̈�LTd�9��AQ-Rm�kC�;��b�|�w;��Խh����,��M�E~���ٳ�P`��gS�~IY-bE*���.��Il���uhn�8W�cP&�lݺ��J��ᳳ����{��,--=	e�:�tqPP��c!EWl��o޼��f�A0���Ǧ1r�R�L��&�������?S�G��5�O� X��III�m��7Ç��9�}�`�S�������G��F����36ZW�\�����ڥNa0T�Er<���K^ꤲ�x:�k�[�q?G8���PQ@Dq�8#7w�xT�$?�mVAT�8�E@T�����C��^�z���mTW�`�!bbb(���AHnÿ�A]q=4tP��U�tt�6��dI�Pₕ�Xq��u�c�LR�Keu�<��Hz���=��H�MBB��:��?&��Y8�aF$�V���ݻ�#���75uu�4�/��j�݆e��V�ɯ]��!A�9���W�� xm��~XI
�J�8�� l��^�Qȉ��[=������Nԯ�N��:�E]�h�����Ne�^	�f�?v.٤��o������&�w�6��wM���;�ĨYH���� �c��V�bT�`����	�O�IYs��v
Ӫ*./Gإ��p�֬��3=�/�~�/xxd��}��@@��"�1�i�U�����6��#�;65��3�Z8�kC�C��H�̤�9*p�~�7!׹�X���3��;9$Ե�g!�B~�RL\<��8�Lޜ��Vܯ��oq�M Pn�|+� ��1�o-�J��/j�r��v��A'� �)P,�Z���QN�-=��
(�K�@�v���6�_��|8�����0�.��z�O�����z9y���D �08~j�?BN��eee�)�I{!!��P�c�6_p$=jw�zwJe� ۉ�UV�$$nhۃ0���
4p�d��&���1���y�%��)����$��V��0)(ꔛ"� ���0����y��ֱ;w��C�W1������]��!�\B�?�DK�cP_�q8JF��0��&<�(s�A	H�����qU��2<{��'%%%�C�_�2�5�΃���Nw��f��]��Cm/�[�(��7���9�ԴV�|��^؈b'J<B �nX@�hn>^߸��A�����4�h�O�}=:�ޕ�O�qm��O���=b7������u�ʃ�B�O���_�X�*���oGFΓ��v��(P�QYU�?8����l�j�%��u!�7��x�-�G��B��נ���~����Є�/a��j�yf&�zoG�.%��6�Z�2�[E&i5ȹA�C���e�q�"��t�]��\~����PW�'#�?
�h�F��+M����=��B���0�L-`m�av>`�p�������^kQH���$�777\j�;�����88�Z4�K"��D�Q�����jh������+�H����;��	tĀ�Jf��k֤�:�w���³�S*Q���B�=x����I����޵��TeX��_DDD|�"��	"(�6k�k�[9��9�1�>=��kzzZ��1��Z�I��O�I?x�g?>'~����I�T�L:�i�-��x �s���>��m�"�4���yV	�P�u��8��1rLt��U.xY_��}:"�N��]�Gq��~�<66V7T?�6?����h�Z�@�;�cǶ���,Nh���`��	
���W;�;�f3�>�����5�-b�#��+�Fb���¥��Qul�I�C�RS,-,�n~[�8�ڝ�6`��|owE^�(qd��y1(z=	�P��[����]�%�}PQ���/�J�px�&�Cx<FNJO���e/�|9(SB,����g]g�D �6��aq0r85� Mb��e����t�;d��}�y4f#^������C��%������]�=�3 �ǈP���t�@���եIe�!��a;3oUH�u�j�,x���tq�sL��:v�^��+;�I�j�Jص]�[ߛ�!]X�{���?d�l �==bY������Z��^T��Di7~�X̫{$��AG:+I��P� z��Q���p\��ʊ���
���#4^[�pwH���e��8���O�M���������]:N��{�.9�i�D��ދ^�qT�$~��Uww�8�S�(������f��P{�vv�FG,��A���������rx�}"�,��-@X����1P��޵,��E��__��9�D��r�aEu�c���GL�ʬ���I�A
Vy��9�x�}��ʪ%�t�?�B�MM���kl	>�� �pB��~�Y��8~i7�&m�����6�jj������Ux��9кT��E�����Y�?qb<\Z6W6��_'�%�իW/W����l�����-�L���n�@uxF�[��:i���q�C_�cVfݥxF	"��S��੿v����v��jDQ໫���÷�Z�lװu?I�@��[�'��K��D�|n�6�������|�<+1W�l���f8�Z�����靐�������W�z7s���b��\[绺�*P��P�7*���G�� ,�R~�sN�[5S�7М�:�ln��)��\�0�9����N�u-�n�O�Ksv�����D�qο��
��{���^�뽆��[�q!��f�5%)1	=%��y��D�Wj!��w�X��;���@}V���z�l����7\8`Y}���Ԣ&�JN���(�~�kg*9m�3	[�*��� 	u%m��dɒ�z�J,L�����
����qc�[�j)z�h6AUE3��M�n�����X�s��L�8Y>��o��t��j���Eu;�%'�-��0����P��$���2���m7Lq���ʭ��l�������f��6����㭾�p�v���+~��%���0��y555�q�(�g�:m �� ==};[-@��7�?O�B���҆��Ĝ��(�1[��0��^������a�oS] y�H�u!�;{����$N��*����������\�mo�p�_7:�H[4���g�� ��;)��ٝ��_G`��R�'I�E��F>}vj?�Iu���w�:J*��zA\3P ���PW�OH�.�ѿ˥�N�]\\:?~�X"�d���c�����}�qF\�f�h����4�t�A8�رc�5�Ø�\�0��}էTƧ�z�I�?��F&2"��6H�$�����2Fߐ�kf����η��s�ţ~o�R�i "e����>#-�䟆��JS������v�����;�x��̟粆��n���pY9�t��!�5%��Ep��`f����<,��p��k��<t���'�$1�^ `b=��NB>f$�w����]ZU�|�7����W���/_�n�˃l ���\�j���2,�B�t��*J�r�9?2���i^YQp�<�m]Jõ+���e.�4Q�/>� �--IP|hj���a�Ď�=j���`U)1ᓒ7�
�>�ef��OM%@��_�P�]x�I�K!GA��c�ⅾ�=��.x����N ��1r���6effƟl��Lf�LLC&sm��F�(}r�3*+��(�L�ε}��U a�R9��ӫ���S�	�!�0��q�w3�y��ap��N�]�-���l?X߸g�:��t58�e����99ڥ��9p�W�S@�Y�a5�FO�������7�d���\\����r�P���!�g!����f!ձ��\�S"��~�Hs��y��o[��)���r�j�T�*voh�@���x�8T��ǧ����ʈA��c���!Kh�_*d  ��RW�y�k��1�q�G@6��X>�y,iKb�X�K�}F^�q�������혶$��G�kO����T*8̗Q�@�+h�ސHS-�KJ�:�3:��*L�;�a�,D n���������>Y��<Hv�f�Q�$���-k�?�٢W��R��Ė�u��VKl�O��ȼ�����߱�������o�[4C[-�.3��q	q}%4�֎�J+<x�Fӆ�#�q����a�{��FG�z��V��w]Y�gO��&���d��F*�*�F`*����C� _VWW������y-Z��}��3^�<�,�o�Q<���m��:�<[��?6U�H��F1��(��(g>���M�?�a1�'����;gTV�Fك�k:�u����i*���ഛ�cZ�yLG�/$�����"(���D�h#+����|KX�JkP���Q��§_�f>�/���r�$�w=��Tú<=f&�� ��"�#e���b�2�7���9`�Z��N#8}5�_/�+Q� ��*]��(��R珧���EA� b-s3�Hd5��:K�25ZUHh"�m\n\87�[(��O��@#��'+-#c�2J�*����4��&��h��w;�J�6ۅ[�����8�bE?��^bo?�,V__�B��r`b�H|��
Ѧy
�.�r�v�_��	盔�Ѯ]�gΝK�뵨j��!7�����j�Rn�ٜ�����	�m'b��v�
$��
�*a���~�=�s��?pE`�d�ܝa��)����@�,)_�nB�YW�)����^)j�����Bא;ɽ�k���	T�`�;�cMN�|��d?�������~7���������h^�Gg\��{y_���E�9p`/��_3��H���|�ʕ��beϋ[�[�j6��4�$����i��ܜ땔�< ͌���~����[|�׎����@�;��̞�k��[�"�!I�727;��� �瘸d
�`Д��4S�KYf+5�r	J7~���FR������s�)'��p�KIK_��3M�=/�>�:�G� �9��tT�҅ǵ�VΌp���&��(�;�zo�K����| (V_�:e�e���P����<���=˰H~�;fʛ"ףt}��L$��>j� 榬�T��C>�X�.?C!_����p��=ē� �AP�����]��u��[�=(��^�^����I��U�i0}C{{��Į?ny����r��6p�7ڲEX���G�F�燗�f�Q-`+Uz&V+�A�@��_Ҫ�WǗ�F �&�'�J<�ZΕ����')Za��Q�PtǛ۲z�{o)d�4E(gtJ�v��l��A�����z��Ӡ�'�����A���1����*��7���;�� ��=��\y_O0�f(M)����Ȑh=��ɀ�xd�
�/�mz�RƧgAX�3@���7�o��+����Y50$T��̒[%sss}���z�k�����"$WB�h���C�?�*��L��m���-9�X���5���g�ŋė67�C{ZB�@];w�1�z��&���|3�6�';;{�]| \ �+@�"�<<6H�+ǃ<s�L��De6X�_?vx�c0�crM�e��Hޱ�[$�LfЫ��U1y��q�<�xx��P�?�%�p��{��PZ�M�"�-�@r���"H/�V�?!�N9<�ַ2�hR�лɟ��Ȩ(sc#���e�,,,��hy�Ѧ?���>�6��;p��7o���/ �Q1��Y�4�Q�^vMsB �|�����V���>�2�|9ȟ��Y.�h{O<�D{$�����=c�Љ&�����b�DM]}�,]�u�w�VUqM�qP��m_�E���W�>\�0�݉�E0�w��{�#��?w��f�R�V�t�������{��jOgX��'j�-������E��Ӊ�mFo+*�V�^M�������1^ T�WP��cp��I}�	5�x������V�Nl\�3j���Iڪ�a S������#Y�%WN?ѐ�V��+����xL��xqw�i��Ҷ����̳��W쫢�icp	S.p�BS�Un��R�|+�U������;jN��s��bP��O}ێ����Y2����ADՂ�o��W�}Ǧ�u�x���Y��>}��X�x�u�_/>�'��m��:E�^���ϟ7�.l����l��]���6��R�Yû��m���۳�6ˀ���E���V���eVN<�W�z���j::b�]��O����6��X�~TW{�`�VSw�[����\�/D��(ơ������V���0K(����辩�a0�#?�Z8?zܯ��u�Pj�q9ާpv'�,�P+T�H�;}��sSS4���#('��^�}��2[�H.�*�999���uo�925ȦبbQh��g&i�u���c��t�P�rZ�{ �
QZm�i���ҥK�Rbf�0jB�������I�@!��B���� �,�6y�&���C�ìƥ@b�S������Q�m�m��se�TN˹�[�J^�zS $����)<ɂ��Z��OL�@��"�v��(\���x�W����LQ//�Gr�����G��[}�#u{�����	%���0��+eV�VMC���D�6#mϑ�8t7�3(��5������@Ͼ��т���55���ۣ���uXJ��U@D֩���{��ϗ��e���t+o��yP�}d���A�����s�%^��'����|�ِ�U��sڮO?,��D/�}l�Zi�o��]�%W/�8��H����~�y��g�"��4[�+�|r�-TM%Mc6��R�TCV<�c��o_w��[��(���t�p�hb+�III�_^}���C#�M����Є�Y�K�#��W�� N�~�yh�<М�ڋZ>y���l �A�� �RA"<�]-�|l���D����&9Sw�\�]�`���d�V�P����щJk�n&�Df���Hw~y��}�V���h�A܈,�T��}�b&�Ҷm>]�&iŊ�9�%)��O�A�t|�*��to4���j����L9��b�6{dnL�ʖJX�z�Q�r�(���B�)���c��Z�ص旾�g�A������uuu��ㆆ�%��wns_�xHBO�>�V��P}pTFFFj��t6�h��������T�ng��r�6/|	�2��?��OYUW��t�3{%�f]�3����o;X�y�����#��b
��-��,�i7�w�!�FÇ����ǟ���"�������r�6@?�W(�p�eS�g��_��f��E�l�=ץ����k�Ww>9���y#Vc��q��J?%�U��8�f%(�������) ��w��Ѵ�W][
u�F�uf�2��g�����ɝ�Y�X٪Q��k'�U��Fe���N�-�B�dl�Z砤�饯ǝ}+��]�7;ɣ��Hfh�J��#Ҷ���a ���|�����o߾����~�#}�X�h�o���I�t.���8�Ѵ�+�	�+���rfpwwwօ��yks��v���j]h)Ե^0x	
�;�u�툐�硧�1���SI����PZ>=ޚ�刎��[�����J$H�����LU��T�m��I,	

RRW��b�"q�=zM��j�7z:j�K:�B�]�EG+�Zf����wF��ɕժԈ�zy�������߹{�=|�LJ��蘻U��w��~���K�j�� ĞL���MUe���ٻ�VA��z�*���9`���k�R�D.�ٌU ��Ρn� ATa�~KOOϕ<����%�\�\����*J;�(�6<�bf�۳�<l�k�gt&ill-�=�68͍!ںT�׀[쾾�+y�c�WY�y���Ŧ�91 ��;I�p��u����~k�z;;��vv_^YqI�*D��v渖�8@�	x�A�<�+�ŋ��� �def2� ��|��o\�B_��s��B~9�6�9�U0"���&����R�JKK�����Lq+�M�-��P�rz���i}o'�:�V��޽{�j~��^�[LRPXX���TU0˪5,��3y1r'�f�=j��/6[�����egn�G�</��F(��wM���4<G�3nh����/ETQB��֭[!s��JX�hhhhET�S�/rr�k�WA�;ja�K�r�q�N�ڕN)`���;��N��$��X@����a���S��{LR�\`�[��'��I�|��r�������^P`���A9�`�N�E�*������=��M%� �@Y�ѥ�C#���Oz=�j� �JKJ��	N3M<<��^`��ÿZf��Õ�%p}��$/o�e�b������~��pFL�V��9��V�"2�x�������<��-���7���QG�slD.�}�c���{�G�`�{c.v)��#Z����	� 3A*��yi�I�ni��'��҇Em�2�e��6�5_-N�dUF� �����N�
[jPɉ�2��$��Px�����oh����Λ��Ȍyyd|P��nP�FG���,ژ$�(�����Q{�V����t��V���!��a1+�z7��t~K���m���0rn�u��8��Ij�ށI}D�A�o����D3�i�y.+?���<��PAk�ï���a��bP�?��}*���nT��n���FP�hm��H��ijgoof�ǂ �,/7@��s���5�Y�11�����5��S�+�=)�Aɲ�,�؛6��BևT��CԖ�~8t�|*��*���w��<o	뀂�6����#���ZZF:o��D)ceuݠ��+�V |]Y�r;$$��퀚���DChe�B�y>�/D�y�����R�4�`�l===�es���S�@�e)"����C�j�&xWy��9�045`k�0(s<YS4�8 D5�ė�.Ng'��{	�.%%��*<��:����+��&ZU!\2d���h�����AZ��WI�1�;�v�f�o��Z�V˯6 �hyO(�zw��:@��a��/��@�q��v+2�[ �CjWv|���iӦO3��Q���1�?8J������:��*Z^t��^D8q��!dɛ7o��w�xf�ޚ���ؘ��j��5Ǫ�!��J����Sn��,_̢�ի�����ѦI 6��e8�}oo�N�Ү-a��t���_��ca�8���	�晱�a������4�}���!A����<��U�Ǳ]]]���y��w��Cy�RqE`����l���36Tg7f����E��l
���&���:  ��ɒ?��2�&�8��!����&۶�d���ا�GS�1��9�L����e��x�H@�u]h����G�N�8�D%��#����.9�v�e>mG|B�Y7<_{Bt��ߒ0�*u����Qq��á��pA�𖰣d��H�C@Q`,Pt���N��h�S�=YN��-$x�V�;��EUf�ΔWuIGb� S�j�F��4��ܒ��]�� ��(U � R�hU͟C[���S��!L��b� ��q��������j4 �N6���7��xt��pE�ޓ���a���C2���J�����n7�<�U���9Z_1�c�����	�PD˜<�-Wn`��g�wP"�8k���O>�jW�h��8��K$�ԏ�߁��sMT��o"���	�$�M���f<�|�\nL�ɱ�b$jNЁ�ˡ�t�9a�ǞT�m�H��i$k~�H�g.��"�4���17n���I6����o>)>�l��͕}��|����x� �ٸ����ɓ1MMM$)��n��|6�t��Q4�D�TA0/�r�'��.Į���_���Cfl�����Ty�A�W~��������0A
P���)�."������"�Vq��h�5����#�\!�����u|Yҏ���j�Wz�]Q�>�8O� �ךʫz�+rk��7���P�t��B^r/#;;{��`�L���S؅��Q��Թ��jXWU�j��{��r����k7�ő8ן��"���&�9��f��N�ɵ�-�[��o��ͨ�NUUH��!1`&�<
c�W�M�$�w���m	nBJ��|}���D��}��7�&�R�b�>DE{zP�/�h:��!����_�Z��"�0��j��7P����c�ջ�ě&j�~�8U�_�;��~�yPґ��J"*�����h^Ӻ�0��@ظCU�HK�s�旹I�I�����>Lz/��F ���X����2(��:	�����@��߼)N4O�Eo�ݸ5��@~d���Y 	�f���w�׶-���G��c �������vm@1{��y���������ܳ+��؇��Xo}���D礏O>�k���ݷ��sM�2_!��T��i���<By낳M:��ও����0�z��Ɔ��`5j�#��
Q��	��m�^�M:@���(�@����h��g�\���K7�) �/�k7߀L���Y�*"��7�rOw/���Q�����=z�TyB����1�oX��L�UW����A##Z�f��9�����G=|�EO��Ɩ��vS���sՄ�g%pi[4�/���G�7w�e�CK�<�ӯD�Gg8
(��*nZ@X{�ӧk�}��\��-��򭪲��s+�ړS*p��J�34�KE��w: a��F�?�a S;~;o��ic?��_<�u0���Eԯ���P?(͛9#,���x�n�V����or|�EDE�5�ֆ�䖏��F	h_R ��C`XYɧϵk�Y�$M��t@/����Zû~�����{m�[,�!��m�UT|heM_VE{qBu�^'h���@{�ln�)-'�-�K!��5=t��ܯ�7;���^VV��rA%tl�U���>E8�<�H܈J�e��r?:�
[C͓(\�/����pՑh�E�cǎ�ŝ�a I?����T�{{�������'x7�����i��"���s�~ϰ����}R0�c Gl�W��a!������tt�[���&�߯�ߺk�44"��)(�����ܝ2!�T�}#��,D��${ X={VZ�7��x�&k�Sc����L}�=y���,��:=��O����_�"�����G"Ztb��\�m�>�>��v��	������!�{řv�mio�!ع���l��n��!��^^������ؽ�1�TT�'G:ϟ;W�ݲ�)�^���~����2�� {���er�~�����a���;O�f�� 1�n��m}���\A[}�^���jD�b5�0�¹h��{AmiF+=f6�21�~���)�����5BY������2ؒ�1$.�#����,����_�:I�^���YR�I{���B"����̽GE�6�~�0o�=8ߐnot^����]n��"H�*V�;\��b�|��)�H��9�"�'z�x�v|������/'��_ru�[������8���F�̇b���S��T(&�K����?��R�r�A�n�H�Y}�/�(�$a��9���4��������[�|D?{�C���q	=���	�{��Hܒ��β,���| G꣥���_*�B�7��⡣�<*��,"hh��ꚱ�Y��@�pf;�ZW�������U�! �%���0�/^Ƥ?4�!c*fz�w���ߎ@�������}
R(�V�j�`Ծ B�	������T8=>�[A���sZ��h��t�^��s�=�D�QȮS��%�T~��t�����lvh ����N9��1n�u������Ӹh}��-3�g:��FۍU��M�.hK�(����KfA��k6m���{�TR�6�up5�����ƢFr�(�(�]'�h��pj�m����h�����bB[,�c�
�9}l�y�_��C��و~� �RA]Ą���ui���?{F�q�tM����;��Ũ+ܶ rm� ����� ��� l��W6SUy�b�\���DZ�Ԑ6p(��d���~N:��0�Ҁ޲!�@f�|�+R�=���A9nbf�긨�T;�,�l����h�
-��"�� �7����K�eP��RQ�8�O�8���%�P)o/�� ��fYk��L݉�*v�`� �����I*��"T	f.s��q^�c9rǒ���+555�ܜn��n��^�z�*Uy7f7?�Rq�J���!m�%PIn�R��U���J��-���Z�I:�]%���ׇ�Z�^���J-��B�,���vK��:դ��Br�X��Y| G��$��&�V�K���
qM.p�]�T�U�����4;���aґv�C�-0X�摦J�!��\�h�D(�F������:Z�0���9w觽x��&r��~��W[�b�o����2�u﬽��t��4���7H3���ٯ����廰��UUؖPƏ���"eCD�*��v���r����e����2x}�/h��.�Cc�aqޕ�GRԚ�8L���s	�dϐ�� ��V�2��IJE][t+����qe%���f���Gϟ??�R�Ә�赳��8z���(�������㼯��@p�S;p;!�^ǬuF�&��˗r�XD�
ѫ W�����]{͑�?ω!<.�*_���I3��͛��O8�"�D����Wo�fgd�}xK�ѿ��F��R�Є�bF9�Gf�NMѪ{Ƕ �u+)>����`�˃kײ賴O��M��A5��1t�
,����!"J���ns�9��ȱk!D?s&)<2�ulBh���+�G�H>k����[3��X���f&G28k��,�e�.���5�7]�te%�$�ț�^�ƾ� /��l����f��u J��1�@!���Rc3Z��X�/�k������h�n(��]%����}��>М+9>�| ���n�FFF��p�W���k��q-�5�����YSW�ìA�b�@��~�Q-777��b�L���\�Rm����&���Bs6*v������9yF,T�P'Uq����O���yN:8��NKk�g�
��lW�G���՘5��E򷬣,������ds[�������0����1��o��u�H�߽��_���̌H�}��{	^/�ι�np��nh�|�������O�P�cA]袣0b�׈م��
V���4�\�~����X�R�P��<��Im��>�N�"���^C�~hh��3��d��W��:�}�x�kjD]��l�;9w����.��@��?c�回�6�Β���Z=������ΤAȠ��TwBu��Y�.���4���q�Gi{� Ru~���H�I��������伯�ܼ�ҝG5�T>�놠�+?�R�]���艶h�$� �G�j�D���40Te_�3&}�o�N%�_!>�Wg��F{���br����K6���}��ᶗ�԰P��U�B��~(��5����'6±�7����!�AE�^e���t�*�j��K@hؿ����F�cd�4��Pd9	|�
a��x}�ا�*� �1��TBOeU���6oMj�O  }��e�S%A4pd�Q�΁t�ݮ�ڥ�EpC�ѿ��ű�5���?{$~s`5�ǐ��c�v�8��:�R�����jjR�{e�n�47��S|��%%y�����^5j���܎F��p����S*Z���[���;��zC��v����*�Le�c�u��iiκ���S�~����wTF�
>=�����D�}O�O����m^\�v���0�3wwE
�����P�Uh��܇׳ڐ���־Ҕn�V�3x��ܷ��g��c��C��4UN?�s���]G.�?��_6��n��`�B�}O 9��qR��V�dR}/*E'Ɛ�J�J�4�����	��<�_�'�f�G~��G�����O�F�m�F �j�Z�&�m
@(X7A�Ъ�l��J���egO��`&�ܜO��!�z�B�ugU4"��h�TV,i��QL2����Ǥ]�}}}jّ�
-�䢢$�=s�cI��%����J�sݛU����J}>v�)��pA�1�y]���I�rJ3=}���=�J6�t��ܓ����3����'�!�%`lz�����D����a���!@���ґ���&��0A��Bp�ÎSo?�f�))��F�� C��{A"0�u�E���P��/��	�Ѵ��׀�| d�|�[�Q񻼊v\j|�Ύ�s��!	��ϲ�P)�N�c0�5K�`�HDP�����|(��s�9c���WN��y%���J�$�����"�*/AD|M�j�w�7j������ݞ����b�L�l6"���:�	�%#Z�����(�0�U�F���0����~]�믐�cц6�^�4 8��J�Y	�b ٝ��F���e��&��X��4	��sKJ�p[/��,�K�v�p��C{�^��� ѽ�G;&cI��ٞ�`Cc㻸x?ת�mnh��BIՄU�J��r�B݌���L�^:A ���c�|�}�x�f��S�����;p_�S������|�q����+��+z{{�~��Zm��R�~�:���˴�C�8�Iq��T��<6��'�_B&�4ѻ #c�i]��0��ћ�g�R�A�R(�X��yK㊐���ʢ@T%Q#������TG��,�M`������F��K������L}� ��bFf�Dϩ��|�ѿ�鞆FN�9�R�H�$�`K>��?Fی@l��#�9d�ƿ�7���=G���Ǐ���������{�5�c@�<��gɂ�htt�$O����<fiIbef7�+��=�i��'ܸ��F x' ��F��ы��_�� �βqla��Z������g5\	�8S���*�;�C��ܹs@{�Z����/ßf�O<�!������@�zL�ihBj,������z���&{�%���|�L�R¾צ�	~� �T�
Ϩ����od�K8w �vA�TY�4k��E��!p[��s'.dc�4�,(�Κ���|VA��/��+;-[�hA+���z�hÓ]����m"��fblg]�D�^� w}�����0��;}a�z��ϳ��qwڑҳ�����!jN�3�PE_��=��k�gG#�b�-���z�kc��WY
_u�����AAA�"5���P��\j-Z\��ڀrЙ��C��/ӆ��m�W~���v�+���b�jh�O�hK�r�Y����V��R	b%_�j>��F��ޔ�~��y�.�<���������Fp�n�h3"w�=���4#bu�U������N4O*D;5�{��x��̓J�����?��}��l��l�*l�
�zH�	�� ��k�r����d|��1�^�tx��%K|�A^u�B�������m>�	���&��
��]�̻�Zlm*������}�ݝ������Ƣ�SR��@kL���%X�M'���/�	2��J_��`��-Մl�ŶV�<n��,�FЂ�S����6��J�W�0"���'~�BnBKW�ᯁ�~����⤻����N��~�X(��w�A�H��@��ƶ@�啖������$��b�T�`ccc(z��5rD9-/�2%99���E�sá<4�]a�h\��m��S�hΒ�lE퀐�����yF�' ��Y����t�N3�9�'""�r�Kx⡄�goo)�~��>f���<KIYq���1��d��c���������+W�`/�'%�]�@\8�y�1���AMӱd� n�قj\��L�� ���YH�����T��7M�362��CVvG]̶��k7��"�(i��~a-=������x��OO�[��0�? ��V�\��MY��C�b����$D��p��8��卙]@���{���t}�{�x��g��B,
�8/��rBv��G��'ћ�t���� �(ĳ���_y#^Keu��qSX�9��;�c��*�h1
e�r�X���#���)�!�j����df�l56~����c?���?��#j���H'���ߤ��P}J�B���Y�VP.v�v��,�1��|t&lEG�ӡY��w!z�Y_�V��;T��i�o���BuXS����ڏ���Q�`�H�=%5U2,�Qo��Bk;򗍛	D'�@�N%����vq�Xj��nVR[{�Gj�a2���(�������ǡ�N����7fـK�߿ע��-5E4ƙ�*�Vnz�Po���x=�3����,�첲2x�-.����eo�R@����2
�+Κ�)����bxr�K:N���ڕ�� �����������mS�{�ҕ�d����Ay,������O�Fu�eg�-��Eo!��\QQ!��e�W�Pg�q�����;-a//��o+Z���xN&7�>�}X ���S̲ɰ����h<ݾ!#�̘�VԈ_��t�{�N����GR�JC}g:0�#.���UmoAס���9�����C�H+)n]����w���&�;v�y���v�G gd��3�ց/��l�������z�n�T�P%��`�'M-�C��@�r�[u���3�Bښ������L�����%�#��cA ����M��\��qIQ)K�JHʾ��5%elQY&k�d�:�V�5{�qJH��K���S�X��${�����t����>ק��4��������y�!��R�m�	�~h��:|���A�rj�S�T^7.����˫M�-���a� �O�2K�"v����7F�t~�D�	^�P}?x�16��!��My�_��,���{(%�!Uy]s����#�������4z��`z��	t|�l�c[1����w�L�u����Q~Փ�"�.`��a�aA�0m�;EZ�^Ye�^2�hy�S`�2��}n;���X��1�����������{@��q@��ՌZ��B�i�J�W�3���yf[�>e�]S{���ֲ�[�ڨHr��In�{><lq��L�e���}<q����,���\A�E�_\!���Ӆ���;�t|��@t�I���_!Q-XC����o�ޤj���^�-
e2����Ѯ�3��$�c˳��͛(�d�e�=��p���iYY���R�;v@͍�d��O�ty��k=�ȶ��>�a��	�cJJ�kݕ�	��O|Eb�������g$��)�W�
c���!�� �Z�x1����א��'9*�;��wB��*� ���	;�s���I5�y���u�6/�m����M�峗��Ⱥ�5�r'555|���e�R��?�Y�^^F&&&Z��NbO��2�V*A����03��e���|��v�LB{�.��j7ev�  �_P��e�9,a���vv��i�t�g�t�������2�&e[�-�pq�������ϟxh��~K�ī"_�8v�������%ܴv�q�}���RS?��|���V����!(�pA]��9�/J@�aԡ����B�'���H
p7������H���P~�KK�TX�lon���?�	��ڋ�����gDq ���m���w~�(�����`]�jWր�nq��^�C�,���T�]�ꏱpǉp�	�.���sߜf���p�Z�]�b7�A$Wj2,rt ��Asm�گ?�]Y�ɇ�����[�tx[����}�P��x����"Cu�
[l��E6�ɌUo��=��,)5�:���
�F$ ���:����Õ#��?s������Q�3ä~�'Z�o�%a�w����^�D��;�-��H6��1)�Z��nD�l�;wP����=<�>�~�W9=�r�I&�����iA��P[p��g]����	��i��3�R�p��E��>ii���Smh��A
~��8����J��SN����}�/¡���5:3sV���и_u��­9��bI��3���+�8���Z9�E��fX)�����;����եw��?����Q���v�}�k�.p��U��)�t{������m>��?�6.�E�'Ϋ1D�y$���2��w�#MM_|��M���!��#OY}�$q��b+���A�"�M膖���e���t~�6�&4��M4�g��U����jx�θ(u�Ν���P\K�ƹb�����h�"��<9[� 8˵�C**�yyyOJ�GG�=�_��5�`��t��<VY��u>��ǌ�v��\oooQ}�<�����<fnm=�1<VYX8˥���xSw�[�n�B �E��=/UT[ۡ���L��������ϒqA�\��@Kծ�]�7�m��Pɡ���Іk���mmzzz��m'�R���-藣��̰�%��߶� �l,��^��G�
���"�%���F�����KݓySQ�˥A^_��yS-ls�@��EQ$
�%@�F��.h����[h�G-E]5�X�uS�m�Q�`�S�1cQ7�;ޯZ�n:r�*;�yG3D���	h�}]ޔc,�1 P��K�ɐ��b����3�<��[m������Q�����.Ղ�/���M78�����ߢ�1�$EG��z�@�@>�f��Ǆ����Nn���X��MCGggۗ/O�9i�Yo��C:����11�(䡽H�E
tq�LL璲˷Q���U_�}�xۇ��m�.0B�����T'�w�0�6�Җ�s����G�kfv�&%m�Li�>w��h�S�����CX�7�!�q���,�O�?rn��I���mm�2qC"��r�/��a�,��ꁯ��5��&31� go�Um<�l�dõ�k�]�r�g�$�d��l���`w�EBh���@��t�u�Gߡ��+Eee��R�u&|��O�5�C�O'���f|AoBd���	ཚ�W+e �j
��ΫNsUT�����3;,g�J�\
������EQ�*hb�cUr�Y%9���}���t�AX����E����׌q����`�|6���+[ގ�_��!�
3]=�I���,��Ȁb��q��Vp;�����J�]f��b�>�AV��|��e�FK�����*�3�C��ki��b��}��qk<詚T����Z������}���`��T$CX�y��b!'/��}��۷3Pڣ+�^���bQט�mѻJ�y6��I�>'''2\#ഭ@�\E���m1�Z�~�j�)��a�8��鐽��'�?ߝ�:=�f X*Z�$Q� 
��:�"e�o��Wm0�R��U�Ob<���~/�@�pCu]� ��#١�+�
f�#�E��D8ޔ����
���@�Q�?**//��xs���V��e+���5i�y�5۷o�����׾}{]jz:�n�ά����Ύ�#fU��:YZO�zj!�`���Ǐgj�ӏ����[TW'��%
Ԫ��ؤ�.��MP�y0j&���R�d2�^ۦ�ΐ�T��	z��E��p�ތlId������p�(�v<&&F�):갾CP�E�r��K״�[�cd�.,�U���� �v�[�N1qS@�<�ua�����+{���g�ѧ���/f%J�2��m�g�%��"D��LLM��d��Ǻ�@���t��>�ˊ��X?��c�@9�"��S,s���|�M�@l�舆K�Ū���� 3��_B�����.���>hd�w���������:w��������i�9t(j+*̅��&{�|�<M.�o��z�e��A�p����;�6��b���V[���dFu�\�̭�,&�jp����S�H���Y 'p�f��o�P�˗�8ݱ��D�P���NL��kuva�P��D"�����e/���D�����N?`�B�i��$�F����8ArQuu����g��9�R�6mz�5�KT'^�3(H����b��;�Ah����>��Jc����t�(����9�qu�ӧO�ǡ�m�0�A���i�%���R� %�/���*��uw'��$g'(܀ܣ�
�M��m����6�$����x�!D��������q����	\ �͛[��a��vӉoA�f]�&�ŀ��,�R(�ѹi�U�u$i�c��OB���Ԉο�~'�rN3����Rca����e0����h��!����Q�ﺈ_C'�=i���>K���w���Έ�K�����L|�����}%K��뎎��?%~�Ӊ�韯=����ǿ��Kv��+���:�op0y&��b:��Z홐�8�K���e^7?��ć�"6?��ުz`��������@��Ʈ"ss�8�F�Ul-s[�*�!���Xyzn�c��09v�)r�U//[�h��C������pH�fT���"�+x�4��C/0�p\�+�nFo^�����^����=�7箩<N|��nu'��)l�V�%�����;QUTZ���	�E:�v�ny� Hft��))�\ܔ7�}�;�W�'�_>�%�<d��ȼn	u��ϟ>_��	~�����Ç�WJ�6g�W����lP�s
��K�켪!�j{�S���Θ�0�h�ߥ�!�S�P_���H�m���3���6u��`M�1�4��[����������a�o+�����s�L����P˲ �ݨsK�v}I���pŜ>�6��c��������n�d�~���w�-CfZ��;���a���������5.-I:Ar�$:jnnT�_6E��4���Ҳ��9�o�:P^��,{���򃈽���7~T�9?/F9;|��^���^�ADz�{�IX�F��6 Xݨ [N<QQQAV�)�����8%� �0 �*U�^>�θ~�r/�n��O�-d����p����btQ����mހ�@�B*	��m�����)c\�w�b"�����TH=XiM{e�t"�x̂n�������� +#��[u�����5�Vch������b�Z��zmDJ =1��e����Ր	�!�"z��@,�<Y�ZFb1��ja�?R�:_Qv��AV�>4�
�'�@�dj�G�b6w�/�2�<��D�UW��׎�i���ީ*<L4>��(�����o5��uT����p����Բ�[_K�$D򖭄�U���<i(��-Snn������l�~�1��J���f��a���o�����)h����P����ȿA�����ā���\�&���ג0C�.(,ܾ�R7�gb=B"\�(�5��=���+��k�6	�-���S?������&sD��_��<)=��*�`�C ���KBo�_�AA�?��*����N����#�u!��S������[��T�L�'񤣏K;�(�߲����C��M�	��-�}�� 8���}�W.H%E��V�v1�"�:��;����W���B��B���O�CU�u�R��
�k�'ؙ({�lw��h�1�Bᶧ�/�Tx_��z���*������7\<���XA�1z�?������dDe��~2B(�{�A�"�
}h��B������E;����~;|���l��!U%%��މS5uլD�w^�fU��j�_/�Y���)�D>�YUC�X s[ ���CQIvySV��
C�z)n:��"tp`����4/Ar�玿w:Rғ���������c�X��Zk��@U��gq�@���{hf��,��E2PΠET�ٲe�ȷo->=-�i��lM��H�F��N�����^���
�.��.�%�~��g~�R�ˍ'����ޓ3nt�t�*��;F���Is�;���W_��A���0ILcZ��AAveh� ju�O��D؋/Z޾��)�}�p�B`��)#i��l7j�LN�\��:A��Z�s�<ٜ�b*<:�d+�V���S�}%���04��H���v}X�s���pV��hL=�� p�3|��� �`$Lʩ������Th�l@D���b:��th�P�'��JN�6c)tS1��^!�ϫ��/ΗO�.����"3s���g�!uV�C���h)���USCƸ�UUФ��c ��K0rX	���o��:S�{(�h�j�g��DFF���u�۽�*�����g��|��Cvn��WV�����g�rc�!���1#\����r|�89�d��˭�y���E���h�
�=b~�WNEf�ޟQ5$� sB�Fn�Ǧg=-mEzh
��E�4C�� �C��I2����*���2���$�yۼ*o��PYع���\��> �����W��D�� ���qC�12��Vr1�����Z�t �;�P �R�Ml���@2�EN!4��~�m6+�-v)�t�G9��3�Hwv1�ؒ�L��2���;��n��!C)�$����7aa��K\�I�S x*'�.mIv���g�c�w��8Q7�0��,�D7�B����������~�"�g�6b���	�@�� Y�td�3e��d��d����5�r]H����f��O���7�\<���y�Һ��I��E`�R��w��E��̦)R`]�l
���в�XK�19���t�.ߩ��$1�D1�p[�SF��I�.�f&X�Oh�'��BF������>�[��C��$�p��|��	fɿ�{zzV���(�]�6D����I�3�r�{I壣�6�ɦ2B��N�-�_�t��+���y�5�Jǥ6��\��H%,9�ə������~ͯ���;]�6�X�^���Ѣq>��e˫��]�M�茞؃ѫ�P
�P�� �j���$� ��Yyk��w�\m�zt8�I�4#�8��.���\�N����I`²�2��>�%k7D]*� ��G+�PK���^��!�pN&S�+��.�'{�_�jlU��L}:3��`�4��ji���1�ӿL*n���)��.f��6(S�G҂����qbFVb|V־��������}Y���U���:�7���-�u1�l�����Z� ӪU�K���}��;1���G0�g�4�,g8���J�g�w�/��o��x�~9&h<MU����G2�YC�.�0�c/ЩW�����!W�f�d4�����cV6ciiia��D��G�8�q�_���䝜��K�F���[� �<�~���+Ҹ͇�dEDK�D��&wM������$E�e0C%H*���_6��^~qg���a��ɛ7o����g�R7���O���Np��1=��f2+�����װ4�3��� NPH 4~�����r ��^��sLC#������k�Hl��w��w�^�j�Ї���a���T�Z�����Q&�n���(��Jd!�cG���.v�A6�ə��j��.��;@K������z��v��ϴ�3��$�j��נ��z�(آ�"Ѳ���u��v|�u7qX�����z�C9݀��T�C��l������ûS�8w�2kim�G9�Q�?,8���Ը۷׹��4���~����:n{�Ϣ�G�jQ<f�����P�`a/�LBC�\�Z೛D�їM�۝�C#b�)̯,����L2Vn�B��WL�� 	���c�����\�_��}j ���l/��[]Y�8�5<s��&�2)�L&b�
����{���~�j���Ӥ߿��y1�o��,��P����71 ��'"[�r(�?/'�r(-uؽ{wnccc(���ʌ����{���{ƼWǰ� S�F��7�ZzY�P��������2t��」fC��"���N��n�l���]����ig��Fՙt��m]{�c�L���n������#k�N�鋯Y+��j�V"��8����:�$�F���w�Kz�%��;̆Xwvv*u,o�a�\)}����un��,�AyÒ	r�:E�gT��zG�*�w��w�d���T�v�؍������&y�P|~���Z�n�?kP`U0�%��1MRlm���^>#��u�����:T���Q��[f�+�r)�I����@�/�H�j�i=>�2���Y�F=�e���g/f��0;���L�8gcK٤9O.0K�O�?���W��4��������5�O��+*z=�� ;�:��������![,C�	J�Z��a��U�h cn���b4��@5@ä9U�۶?�k���Z���`�+��5O�jTx�L��^�;�w1�}�=N���t595��;�oJ��ttj�-�k��9�[�i�����w!.L��s�Z�v�~��Xj�ܠ���%��s)>�T,T����R%��I���4�Β�zex�K����R
E*B�)_����XC:�A�׈d�7#�e�۷�y|Y�,���ˌ�Dh.�n7SSK��܄�MM��=�٦�e��p�1�BDӥs����~.�	���$=̓���gD�ӵ�*[����^e�xN���]n��B�6��en�ii	�3F�����������JTgo`xY��;"Ld����-,-S;w�Z�FJ��������~~�.���T{u������1εp2�3)��2����3�l�'��e}��뎨��WCy@�-��w#w��.+^F^>��!PVY����eo��0wH�G���u����s��r�"�
�.//�È��~1�$z�μ�>��s��1�<���i���M^EnAU��D<�?��eww��
�h��z_�8�##'��2>��%F-������fl�UÜc�l�̗�f��2�KAsV��I��ܓ<w��6sKK���44}1Z;������322�[�[�tA�]��^�f�iF.W�5�:V��w3:;L.*.ދm _�x���= �\�*7����O4��N�� ɝ���Y��q���][�� #�<������K���σ�ysG�s[V��r�?�q6�ĸq��H�<���_��N��-7��)jY��>׫��= `b����� z@}y�� ����m�f{��Rpx�T�E{��P�MR�U%�#�F0�L��/)�sHEC���\Y�V�I�Nk�t�L��d�i�Y�kgM����~:��B
��)��8��ɛ���PH%��;��SߜS�ֿ����	��	5?�S,p�$7�8nѻ���	I�h�F�Of����1)t��kҰ��N�9���k�T���<��K2�n��h*ıu�ge�޻��v*~[s!��Ȼ��E���:�:ׄ��G�!��H_�rAlll�AL����j͓�e��(Š�A�c����EO�m\����4��)�uܸ�g�;��>Hs�*#f;_��N'ϜKv���3��/�x|M��p�ܗ�M��
�k�����ѤĔ��������Wp΁h6�R��ك\_	Dd��q���W���j�R�i��0��"
�l5��|q8��{n�����}��͓G�����䍻'��ů���u��y���������CZ���(}QJ�R�V�O���9�����ﳐ���Ѵ	C��.��Oh�v%(p��"Hq�
����zV��$VV�5�CA�v�,$�7���:�����Ѵ�ꁣ������,?+�'��P�r�����WY���@���/�Fv��27�L���j��v�c;3R�Iz@��|==��c��а㪟���ˏ����8���¿E2����܄�q{�X����a��΢߿~��X0�`O�)H�K��~�ɝX,#�h?�V����L�mN@���p؁=����v�v�T�4c�����!2�,���X��+c�[�Pn��G���|?�Z/��t����8:9��tP޴��h��
z�6g����'(E/&@��b(sh ��FmY��mMn=��#ﮔ���pɿ�k-s�2�0�{5 �2D�=٣K����	��M���Y�Td�̖\�a�hr��=ep�ر�G���~LM����{�����l�`� �y����	"r�N|?�Y�8��c��/#�$W*�_�m�;=��S���$�ʹ?��ў@��k����P|r$�$���KHEI��<.!�o�W�ou4(��\"��U�/
��WR V;88ܦ�)cL-;F�F�n��^4/���(f���X6���������4\�rhF�$��@��n:�o|�`��+�Ru�ik�㍟f��G6�"�fbz�k*�����i�B�Ą��hHk���^Eee�J��(hh�����x���Ȼ��f�[u��B�����>he��{�wl�ؚ�'�Yņ���^0 �Bj�)��m���Q�2//#4r�a�ӕ즫N#���!~���M��˿�KP2�<�B��Jݣ�t�K�� �����f[S~߮d��� v�X��K�y�#�=��}��D��{���"��/��M*)�J��v	���Ivv'(�",�7lk^�_�N��J&�>�Z��$��_Q�bA�I�W�l�W��x������U����u��u�&W����.Ɖ_�Q9v��0�ˡ�O4CZ���X�߶��\�ꁗ�.�"�)��yɅ��us(�o�fԝϻ��k�cUS�
z��1�f�$5�==/uo����	����v�}|<+�ͪ9R�O���[Y[�k��f됈�N ��VV�?<�p
����27��'7&��.�����δM�z=9l&�(��x�c��'����Z�Nn����0i���ׯ�$�#s1��o2�{�MG��0�P��S�G�����|l+ҋ���E�8 2�ӟ̑��5�u�32K� �]
�mHI�źs}r�W�0T�ռ�I�C׼&�qh�8;[�cz:���t�l�^n\�67[����oh�d��"�!N��@���_]8���&�����T$*��a�BX�8V���,��B��Y�X;������Z�6�5n�m����E/���pwW�	��$�m��{mw04y����K$6^����M[����w��fB��P�,��q�4'Ԥi�U�Do�>p��v���P��~273��Sxߡ��ο��+P�9����!uUh��!`6D���?��~Y�q�h�F*Q��Ka���ɐ\e�ph??�h���}�8�y�8@�da��G
����0�}Q�3�S'T%����D��ʢ~�|b!PG3�#�?/i�B�@���h�fy�%j����
$˴?��h[�ǩ��FT#ğ>KnG%����-��X��S$Y�^���+Ի��P�L4�=@6G3��� FP��2{X�U}hǿ�����)�3�j˟�"݅�h7���ssGA���<�*�OQ҉W���^�STX��9E����T'����<��ğ�0i���6j����������9�'S��QZ>/��� �9p��)�	D��!�ݜS#ny�W�u��0�fI �5{	�����<�wt`]M$ذ��lܡ��A�� H��a�����c1��P����_��d"��ı֟?Kn�J -����^ԍ�"j����	�ի�U�#�q��1C�>T��o�����SiQ��G}s��x� $q�RX,cw �1�mL��������3k�����#{�AԎ%G+Ŭ6�ѭ�Q���+��1l�"����m��(gS���Ő��l�ǎ��N=2�}����^~�'uN�@�رT@�	�h1��Qh�tmva�Y-��=whz{����L�(6j��i��q舽Um��2{���Lc���t�.F}j����؏��
P#s!�_�B�|�F��_�:R��r:,���[�Ti������i�dkk�	q�tү��J�N`j�8'j��SF��^�S튜�S��c�@���p	3D�"�h�R�m� �5'±����v	��2��W�`ћ���H�Ygg����h��$/y����z��R�[��;�@4\�������4^�yq�;�Q�Բt�K�2q��ܛ��]�v��]�t!?:�p���-��y)��U��M`}��i�%K�����ݵ��1%�����u����h�>al��cć&cz}�f�p�I	��:�W/���������e;���c�D��l��JC���Qޭ=)p�n��9�>-�yT;�/�2�R6)nķ,�ŧx���Z�_3��RF|ts��������z�i��`issū�Z�(t(%b���^UYƒ�2����wg�
Qw*T�v���[ڳ�<y�dr�WuC
�m�-	��� �Ӛ�R7�
�2feeV�v̰:�I�T'76����B3T�g���\��c�������-y$Î�yh�XX[�Ƌ��2KB�i*t���p0O�*�.��%͝u�~q_bo�u������q�CC�d������u[�.s���1A��o+�`����xm��`IEE�l�L�c�$�J����W����O�x&�b�����?M�N�׉�*�J���3��G��e������k��Y�LF�D��̦D�>��]���%=�Iae��[1�*�<������@�ȥ�!Z������� x ؾ>��E{�Ņ��8I��:>=Nqx���`�)�q=xvM�e�e2y��>O��L������?�*�j+�E���Uy]Cпx�d�e:zkH4�yì ��nqY�C��R$
���^�݁I9��6mB��N��u�B9���&]�3뼔q,^��ʹ.�"�yX)f�jo�s����q�&y������?+����xF�*�@�(��
�f�̬��ē�Ca]��?����CS+�S�AN�N��~)�#f8�|�'lq7�\Df���e����Ɩ"ֲWJEz�Z��Q�`3l����#����ₜ܇&�U(��B���<��D$���_ȩ�����fY_�r�B����P7
� D�
%�}����h���Qh��OFȯo������LLLF>��|Q���P�y�qvѯ�-�:g�2���;TQ���U�3K��)���XV�.[o�T���U���w�6Z���5ۿ�m���b��`ͯ��G�Ï�f����#�Fխ�W�	�}x]�$(k�dDgg:�����`3k�V�WA�=��_5��;8��/��A���`��кF���s��X�y9��x�M�ё��-A�5��ZA��
-J�ȵx=�oK4V��R����^+�}�e�i��hz�����މ�j;nO]�xq8z*"\�_a!��AN{��Ƹ��Q|o{�����`q;����%7	x�܋�tz��!1IX�6�f�}���$S�8@N���=��i�S��V.��Pq_���:H�۷���O@:%--msjr߂Eq�8~TQ����4d����Gp��C����x��S��j�<jҩ�C9Z� ������/�����o~�q�� m�O�4E���Єk9T��/�[�~�s��?f�T��r��W�{��&]l�@{&q0o����2�u���Aǫ~��q���w�'���VWW#�@��Z4k�۱��A�-�F>��0�
 (����_���q�Lڗ���Ek������+���E�F��GWC�d��"�xrD����4�����ѻ�E`i�̊c1�U5�J�xJqF�E�1������g>�(�'�^]���_�.�yR��bc��MOT�YL�,�(�S���/��]�P?���m�h����k���
�����v�9�2ơ���������
�z+Kѻ����8���>�i���yr����2?KB��v_q��մ� ��I��i��YvM00ff�A�ir�����3��z4���5���lİQ� (���*�Fjݼ�6f����4>�T|�=ʥ=�ekd�J3x�U��hc��mf��']dS��!��4,���ۮ
���z�N�y\���yU祜O���h?�W����i�h�eX\��8���zl�+�:b�ò��fQ���� �WVJ.��0�\�jolE���Xl�js�R�ǂ��+>�Si��1�bu�k!'��߾M�=�d9���G���MvF�ˢ>�R^N�
��Ц��jҾ����qwr��}�(	�Cǖ?^�eH\Qln�T���x�&���ݽmv���0�S�+=���v����v?�Х�I�#c շGX�/5X��5��iXXE�0���@�v 2vii�N@1?K����(4���x��K�o
?�����KQ��zҤR����2�|�ӆO���Щn�O����J�����.���ؚ.j��P���}B�>_��X���g��?�qddd|�(�Vu��:��8�dT=����m\\��,,>��[z��[��v�MSd9��\,y_�ް �S���1h��g�Zs�8�˱M����6pT�=�;H���V {��O�"�ɿD ��yu�6����?���]$�����B�r�:͗;e��z��b$PS�5����w{hu%��6��i��X�k���<�X���U�(�q_D�/U���8I@�Ᏽ�r�޵�����紹�{�M���J�E�����:��Xj{}ɚ�c��GS��χO�=�=闞�����k"��?��@H��T��Y���q�mW�T����y�U
-���Qnl��l�ws#�
p���.v�tJ�c��!���IF���۟$�y6����M�L\�|��Ea�9�k� l3���f?
i�������Q���y*�R���7����R暵Y���� �i4u�կ3s�fɿ�|̴�ᩰ��:��ֱ��k�lͤ�ß�� #�k�V�=+1�0��q]��~V�r*j߉��7���ky3�ZZT�$%%�HNHs�=Z�'� K���'��)��z{��с�D�w�=��R�!z�����Fv��+�W��ʐ�:�e�ն�vJJ���x\�k�u"��'p���+\�+����(�aԳ����+�T��F���b���0z�Ə8��"V:
���n��C���l'�5,����	})
J��̖G[�6#vs��3�%8b������v��!$�2M7�˼����X�2t�ʾ�&�ڸ&-�!�k>���wa��
�(b�
V���6
K�.n!�<p�Nz�3	���i~�{�́}J<4�6d�ӑ�V{�P�_�<5�J`-�=��5�ɜ�_�<ئ�.��|���m�x�W��DB���99�X�&Y/O�!���.	z��~w(��`F�pZ�QØ����J^"��p�'���q��Gr��P񞆒�����_ߨ�|xN�?�X7��B������G�3nd��傪�v]E��pӧ;����/�i1�`f@y������k�D� �%��~;�̟Xy�#�L�)���!oQڷZ� û�S�{��ԉ������YVH��{x���s���%�� Ԗ�<�t{�M�3l٫y�`�1�ϩ�������޿��H\1��H��Oַv��K߹s���I\I]=��;�!��y��,��G���P�jfww�F^bD�
;��[��h��c�፟�7�8����II��ҥx}!� �a���������= E{s�Gع����!�%�U�p$(��ӵV��C\Az�6n(g����7�z��	�FNTa4�UO�m��:�ې}��7_�^�*m��y�9vߞ@H�=p�L�:�<vѣ�sɑ3�=���A���/��Ï9��QF���y ���g�G5,?����7笄D���f-�
���J��M͟���]	)6�߁f9E��(z�0�����Ĳ�����ӎ�~�)�������w�$�l�Z�n���*��G.��g�& M0�H���N��Ț�i�\~[�|Xē]+�  ����.z[���E�*� �����2ν�� ����֒�a��L�Z��B�2�
��@񱘽��A� O�X�y0����.t����v7��f����س<-�.�bB�wԶxʱM���G�\pY&�{�o�"k����ܼ.�:��v����}�p��u�3f�'^9�ץ�C��{�ee�����Ž�mjkvb�k#z�)���!V�M�a�z�@��0���g�gO	� >}�$�̄X�v�m�Y=8t�M���)�H���ʒ�բ�R�i@W�L������N�����3��i a�p�خ�$���v�yS�a���g�V�$Nr�+/w��=��N�5��m�B���+�B��O=N�yK�y��(L�K�M�/sB������a�++u���er�p۪<	oX��L��z�M��p��vXT�]�^�6G�~}0h����s�]�����>�ǌ�_��.�Vi4f�Z_��1�
��9n�-wb��錃���))2���ucܗ�
1��@�4y	2=H��G6�gp
���i	��7^glkw
���3��NV�n���ʤ�u�B�K��N����9Z#���g�KT�"��Pf)���A7Aޯ�=ASR��^`Y�M?L	0g��;|l�?�]x�`P��<�s�O$ ��gĀp�5]�e��`��ڼ~m�А"����E��#+}d�����ǘQ�z%��P\��r�U#L俕��bz���0D��/|�Ty
�}����������g&���f��S�+9��n���;اq�F85�Z�j�q:!Z����1�9��Z�;����{����6�Np$%ef�./wz��|�g})(����Щ e��=�`�G�v�����	3>N�f��^ġD����T�3T4�_�Rk� ��I_�զwt��"�?q(�:㌪P
A'� ��E�lS��z=��2i�k����a��P�
�y��!�^��PYw�Nj�bt���􎩩��@[b���e^�2�A��@�u3ͻ<�%�i��nLa'@0��������a���g(�`<	�.�o��:���d�׳�u$���4s��u�ͨ1s��T�:���ݻ{�F��;������>o�|��(�I�i�:EhYo�k������jo��p���z�4�a9��G���׎�z~L�5䍢*�6�?��X��a��m�uu���O�e�3h�0ve�M"+����:��>MSg��5x:�]��v!��{�n�x�����W�Tp�xlJ)�q�m��S��L)����wC�F +}��+�f���
�wh���s�k��9��`�6F��;(��.n#��=����C�	������`�j_�l0��:ES��h,$<�~�N#f��g�j��p0�+��O�T��c�e�nA��!F`�)r��l��Oc������{��ۋ^��^�8����KfFu����r���wy�v�e^�e�]R���(4|�m�E�ѷ��A5d��!9_z"X������X�y����ʓ��d/-�B3= &]�N�雯�}�n@�'���`QFTߩ[�Np�{�4 L��WL*��{���yrr�XJZ����Z���D��c���R��`b��W�'�?{.I�����7�~�ʉd��^��=5ϋ�Bn����x,?��m*@������M*5sqP�ʤ��a{0����S^y=�j�%�/�E���1V�տ�س���W�^]O-$�c��ߓЊ�x��q��<�ÿ��6�EH���+��r����I�sR\�����0�[c����N��ŋ|��{�j,�d,Ve!Wܭ�	B䈓T��c��w��o!
Zs�gE<O��T˔� ֓Sޙ�e%�i*�لvn��ǓiF������ r���䞗�at-�z	'9A��!��Ke9.ԡ׬<�A��wU���A��s7��V(C�+�Ǡ�%��OF�r�*��83Ѽ�H��XV�� N?WC��"U9	Ĳ�t�G�K��q�"-H3���s���E5�6���OB�SRR�	��ΐ��G{>  ��-6�=�Ù��Bm�Xz���z0fk�� �q����r�j�6��r�v< �2����Z�w�>@�b�WВ�侣a�R� �gFߦ�:��:%�5tz����|_��.,���K�F-�������i1�#33�"�d��-˿@���+�+�k��_g�}�_iW�sG��f+�v̿b6-�.��r[�S٦��ZAM��}L�(��6e����YJr��z�S��� A�����X)��먠��J]�cG���S}7�_��ŀ���T�!��������=ZV���ݱSSO�5h�Th��U�3�ÿZ��BM�f�N���������G�m��ۏӶ���;�n���7��&��+�P�Y<�f�B��N�����p:��<Bz���w�\Ȼ݃�9׃9I]a�T�)�-�0p���|+����+Z���D�QNV���}�?��#���te�u�A��g�,]�����p�`T��v�keت�~H��|�
65̮;@�:��g����zy����0B���V��Yˑϻ��O�k�<iwt��+�/3��חL�hٛd&st�E}����~<Pb���%%ig���t}��!���X�9��Rh��"ע���
��ChWy�����e;]�����nՔTzhw�֊�2^1�3�zj|ff��Ӂ�Y�����r)_�<�t,V�P��[�,Xj�qܘ-��TZ	�y��Ӝ��@�� �"���%P���>l����T��{�����z���+����Ӧ�gh���/Z<w�F������r]�Ph�=��b�U�zX����wƊ�N;ǣ��^�{%|4���s	�!�l
z*�� ,22��!�$�(�̖�_��%r�N�Aʿҍ8b����;�����5J������7ꧩ�NB�Hr�=8����Q��j<�ֿD[�,�C�,�u�6����./��D�:�UV��� �V��=���h�"V�����3�-�r�mA���h%HI4�	�����߅�3з���I�}tg��A+4������]�{�MCw��;�&��@�����S3[�O���W+eT=�����#���Z`��� ��V��a/4ڨyT����}h��2:�h��3:�m*a��ևV�}�q�F>��?�UQ�KN�f2�]�a�����{��֦h�ń=��J_��/��ս����$M�����N�J����\dP��<��������9���w'����h����<�W����3B�uXZx�c���2�m�Rr�~C����<,����ٗ��� �w��/��^*Y��e��8`�=-��n$���r��q�y��(g�� ��q��L:�����ۨY۳�A����Ʒ��y�k^��s��P��/~�>O�Ĵ�T����T�S�(y���En���>��xjy��nQ��h�5�� ,�KjF�$��'�!yڰ��P�*O=�79<�u���X%���@n6�{٦���UD�4Zx�C�����ا����_�<�u2b�ݯzh��+���3�Ә��Dz�1�s����ron���;����n�o�=��W[Q�l;??_{�Xǈ��7�	n�jZ��h��ڶ�T�P����6�=1þG_�u�"XY�l�`0z�!�������OwA�z�?&�:��2'_���b*�*�*�ga�zz��������"x\��H�I������cU���K]�͡8]*�!�|;�B5v�gp�2�3�nn����Qu%�Tnm{k�����J�)�H�
!�2g�<�SH(2e:%9��y�2%ӑ��<��M���w����u}_�*{�k=����������y��� �M��~���3L#��8�Gh�Ժ�^>u0��hyrU�W6ve����Lh�ڧ΋�2���$h���d���ƶ��F��y�V �.��XO�{L����y��������v������o�3D^y��{&�ڐݝ|D�7.�����?�{z�w��w��H���{��|�����4v�=��;���6+�S
��/�(�v���Q>��N*�2do_�7�O��REj;�g{��R�{:���nn������u �~܋��B��L�N���)ʹ�߿ӊ@=�[3_Ih@��czz�����6�j� �ȿ����x<EYl'n�3�n��8����|��J�ӣ��G��U���s7so%��X����@
�_-Y��c',������D�:��ܡ"MO�N���UCv�������8�%]��$zN�fS�M��0���:�8���q-����n���~_;ww��65���~_&JԶ��z[6>� ����?��M�*�K�&����D�Md��L�Ulkn?�k�Q*{ӌ���i�{��x���{'i��)y]�HZ��b���ʱ$���G�~;��l��:@�;;��5ǘ�d"�� �2۾(�̰A� 4_n��*�>i�{�e�<���.V���KS�c��I�����"V�=<�G��LĮ���ԇk��DT�����@f#���k��Ag��x��aMu�^�ou�E���qt`�O����=�=��:/E�����~sx��P��yapԗͨF��`c֧x��?F'x�>ǿln����g)�\([�~z�馨����-�LL'^G�x�+��{+ȯ�]��.�z4��,�]|gI��H؏#�AD)�u��-<�凩a��w���8P#�C�p,���|�p%�!޸@;!7V����.�T�ǡҝ<��_�%��z�/��j�'n�:�K�c�G	��gc�_�0�u�4�]xŹy�C����[s����Sz�Oz��%N#���#��G�W=�|�*���^t-���=f�s��(��`f����/�{�����(w��Vδ`hM�'xC\�ja>{n�nW'� B���=�7��J/Ǿ�a��&߲?E�c�������V)���5��KY&�Uӎ�#�gy����EK���^��xL����sT�Ǔ=��E��ru���DP��)m#��f�#F�	=�����i����%y(g*x�o\<`j��j���F���F!�+��>����d>
�f��
}#�Ī�������E^����\.�a�980H=C�P�=zf�%po=�D������G�mvڄ�f��ٲ��!Ҥ�ݝ	<�U���~��2�0�%3����L��d�wk�^n�炷��
��9����z(O������ �����{�K7D�V��[o��s���/+�U�����P�u[	o�X��m�#�-5d�%�yz�,5Vi#PE&�M.���f�**|"��E�"��3t�����o<L���pX]i	�Gɀ��F�×��|��|���</�P�FJS�R���G��?�Pz���kl����޻�{����kY�@ݏK�� ��Qij�CK�3��%R!��w����,=�ZYɃ�$ɓ�۷@CDL�~�[�pt�b[����)m3v��o|�Z9Ϻ�7��������踙[Z�r���@E���2��{�k��Eh��z�V�]C���PWgJ�6��[Vw6��E>��8sP�P���h�	�x��[*�O��v�cc��z'S��@���Vs��~:�@�5u��'Yrx�拨��l�_��?�ڽ�nq��("L؉qV�m� ��{�(x�2��c��N�����6��ǻ:G~���?O[`\�����]��7������T͔��)���8�m�Q��(
ն�,G�s�Y�R�A/��p�FaR|��p'����;��٨��{`ew'M���&c�u������e %�ݍ88Л���r�x��)��������G�]��4|��,:d�zRh@iK�ݍ]��c.q$#1�Nr��as�d�fJ�v��Xo�h3�)l��Eb����q��B�_S�]]#��S�����#_���E�����	0Ϳ'n�4Yꋡ�����ϰ�FOj�o����W��8�4۪k�is(���7YH�v�e�?a1ů�R��+o1��<����Y �{---�}}Ǣ��8�TN 8^ZG�ot�I�	�����g��0���M26���24��I�K�h���g�t��P��)�Q���Dﬞr\���or8��5��F�l�j�9^��y1�k�=&)Rn�z�hʶ�ҏZ7��(*�y���"Q�}H�'�2�/�I�DI��y��6�=�Ex��9�C���QZd�qzl�MFq3�t��-c�E���)9�hn��6��*�-7���j���'��I��
(/Q}*V�����,�8�����""D
^�����%}�ZdV�%��5/�J�T���ÄV��*�	�ҔgMMM^,�bt[�� ���L��CHՠ������V�@n��2��Bw�<����
N(��X<|O�9.����Sa*���|2뒀����thۑpYa���8����:��tN�XZ^�$�Dע�!67]�h�*d2�X��5�-�{��QG$͖
��7�3�uD#�`��p�9Ξy��'��@{[[++k�쬈В� c�r���g���l��X�����i��ƥB
n�1����Li+-��8�(Q����-N�CC0(gi�f=�1A`���Ĕ���F-�{z�}D v ��a�m�� �LK����fs%��=��h���*�W�������Ъ�y�t�r��`�1ћN�}�fe=AD�m��Ԗ	$�+E꿃+���
QI䂹|�� !�>�|:7m�]̺{M��$�aU՛�v���z��[�9RI��ݝ�s��uw������/e�����������b�p<���J�)��" �|��φ7P���<U�ځm�������,7�!q�/#m�Y+�-$����rk}�n�ĩ�����?�t;|8����. d�	ֶHl�H�v"3#�~Jӧ��fvu���O�����Ig#��4�ݪ�N�j�g�Тk�[�L3	�� �8����Nqq�}���(c\n�����잨!��:���h�}�d�O�#��ш�d@^]�q2�U�y�0=9���kL뉟_� ���qn��ǺWw|��N�C�>hV���Y%�+�ɼ	�h���>+����p>�:�R����jѝ�A�|�^���bIv�,=�ZL[���~�z��W9/��p���	��B����T������?{��� � ;n�n{0�y�F�&L>�QDvm��҄8A?�*[�̗6��������Uc�5؏"6-:�-���V�I*�G']�AV�8�G�;=;�Oo��zf��y�P�N�q��6���������v��4���$C�v��3*ɏ��af�#_�V����k���2Q����_V�)�QNJE��GB����;F�L��4�ۙ������nݕ���FC�g/����r"v�k��l���39�����S�ȯ�����q]��g ����e[ngh߂b�NbH�d|�A���S�U�'"g*��#�.�#�����lO�:��y�=3/�#���.�41ISK�Kp�"�O�1L��m%��F����(>Z�9���E�NNN�<��|��ѵ� <��!W��̨{	���;�V����	�t���*�s]�8����r"�z�n�}+6����	��`$[����S���W�����%?�_sA�Ho�+{�R\��tZ�˖1n$�<�����π)�U�#�����@:��ȁ�j�cu��Һɷ,s�����Cј�])��I�lT�Z�9F�s��N3�P~~��9~��⁵�L�L~�=YU�)� ����?w����Δpխ��	1�"vB�!���������O��r1�:v�1�#�Gښ)�H�NO�lc|@�d�ܯE��g���K�"���A\-� ��Skto��g<��^�}����|��/sVZ��g�߿�����fV�V����ąȩ���������_c�N3d�	v\���L��Pі4��ΠS�t+�Q���#�3~|�Գq���uAn�$�f�:w�vJSHl,{fnn��S����S���eh��h�^�M2;�^�OhLr��hw������>e1gSs�T���=4����Z�F���7�г�9�inZ���i+yhL·�+2����I���
��lX��م�s���w��)��R��H|����p�ʂ��S@���z��gH��^�W2۾�6p��Gi������CA��κu�N*�ܭQe,g/	2���4ƥ�f��o�Ϲb'a��@Z.�8��N�/
�4P�W��9�illl_Iɓ�&�����$�NJ��'�����/
./,�Q�;As'5f����uX��t��I�/7l|��y�*��qB�C���(���񔮔<�&U9��U��t�y�vᲛ��eYjn%)&�ra�	��v�fP���!o��W�O�m�f~.��~���8��I����m�����)���z���C�:W#25���$Xe0c��D�����Pw��D��������gZ�Q�l9=�}&����w,��V��5o%�b���n���e�<Y5�?ZQ5dR%=�a��zN=��+ �GM��=����Q���sn�ٷ3\�=6yH�Sx��s��h���d�.�F�ß��a[�fI�x�Szݍꨠܻ���1sHռi��ƴ�S��]-(�A;	�4p��g�Ϳ6���my~�L�Ӄ� ��|ȗ��ӖO�%L�ݽꡯ ��C��>(���y&j�5���Zzh���FK�^���zMII���^�e��e:���7�98>)&�SS<�����XQ�&1P��w`�	C�*��L��$DHd���k�tήT<�"c	IS�6tus�!O�]���EM��ots{"Qot*8�u�n���tW���8����9l4���Gw}�LI6��Ie�\�7ꇘ��)'5�z ��|=D�����>]jp\2��+��4���>��t�ʟ~���*t�{��
������}#�3�d
�Q��lPV��V)�:�-�S�M����-��U��_��o7f��|9�f�9�,MJ%�R�l�/���rb�&�xv�T��Pe]�CHf���z�)����]n爾�P��C����I�(��(�"���"dK��Yr�W\�gf�7M8�&�Bȼד�DJX�z.�·���z�<����e;ry*J��L�f�i;�4�so��fi�9���a���hW��ӕ��ŉ��+G@+8���1��f	��%��WGM�J���s�?�	ypF"�kw��1y*ͽ���ٶi�k|'�,�A�a�����m�-51'�KD�ڍ �ʏ�Γ�؁����L^����k���0���.�7pi�q������d(��>{ۮ�#�~l�t; ��xh�P(m��q��+��Y@P��#0'�p�>�%�5�f-h�:���+쉨�>�4�X"E,8�\c���\f?NA�z#N��o�Ҡuwpv�<\��I�C����ױ�{�Bs�h6��o��e��C��ɷ�G���ft[V��:��E
�oQZh�w��F�S�[
��#b8c&�{����Z��S��Aw+�.|@�P�]j�[dAV\� �y?��GZ�S����&�ZQ�x>��3D��U�=��=�� �����j2����>p9Z%�\��p0�<K#��S!eeb�;&�AU�s@�rk�ro������_*i���o�i/�[�C�S��n�kY��݆�	R���=�-�H�>b��"[�n��Z�T��.ۚn���&4ƣڪs����C����z\��Et__l+�z�Ll�w1P�PE ����޻o�@82 �EK�@� 57��M��]<p�P���n��c�ج#��<��� Z��2|�Z3�\P[ppp9i�K����hh]��@/r'Nw�wJ�x��A�����h%쐩�)v��pK�� �*��gf_��f:]�{!ߚAj��gW0�X a}2�L����=-�)����������d�k�_i>���};���u"���ENNfx���d�A,���Q���ޜ�u^�@OdL���g�F>R�<���s�ι:)�1�F1ei:76\�^>pa��Gwqt��훯%�e��&�n8	��Q/��awF>���w�k���r�

��C��a�ٖ��膔��v�$�t�aF|��Ds����tg��˘�Nn�Ԑ�6HCg�_���In?�s	��L\�H�D �r�ne����k�+..P:�R�ۤz�x��_((��h'��Kl�eb�]TP�L�
����+X�S�Z�W/8J��:uA��V6�\$d��Sk��x�5Q#�/(�-]\���:J������L�!^-�0ǟ�
�v�|F�,I�i��v���⪍8��@�3Q5��NwŠv�M�f�1��9�V�R���� �~i�ɹ��YU)G�u�n�U�uvg�_E��tS��"O�w̥a�f"�PK:Zu�L�` ���^��Ք&�Itg���o�'��%B��Nkc7(n� {tq��V�o��8u �\��w���.����S���O��u0C���&Sg[�5���o}��p�Q��!�]�6�B��kS�;���S����\W��%����񬉉�tA��7�d�z��O�Z-�Ln).rG�I��BTO��^�SI��9n�/z1�k�(�M75���;�>��q�G�`ZV�9���^m;t���N���Jc|��y�%q��M��ih����*�b�7:I�{��|40@��Q#�g�
v�?��$`-���5�ӠI�{��&	��n����V�>��5P؃�0��0aƨ�3@CYHbb"�'}I�=�<��WC��pF�����.9C���tcA�}.N-�|^����>�		��lb��rv�	c%��3L痥oH�jvU�6�}��i�+�kǨ��l��O,�Go���>JCx<���8���g��ɼl:�z@7{��g��o����9Ҡ�+�Ɉ߫s>��aI��(yϴg{��}\���I'���N�ԋ�c���N�>��B��h����	�5̈ܬal���zt�����n�����j^�:![�$�.����l�����������ch��)m�b�I���Xkʰ5�1�����E��A��^Bb�o��|��B��y��&];2��|<P��9�}�N
��0?��;2�������8Փ�� ��� ��%������U��O����e����i�=?b4��\���^�S�=���<v�3��kf�\����JbTvS�v���T<��� c*^"������r�$��-`�u��K�+13��k߱@�� ́T@�$c�\�(mMS=�-WOmϳ�גϣ�$&1f�A��?��ްtT�e~�x+:.>�4�a��,7|}�g�JCڄ�!�%#��Hbr��
��U+�r}�G@9Gǂ�4� xm�h���:���̌�������}��Q����Vm�Y]3yX����3�X���|�}{^��\MILm	[ݾ��5%zn�i�o��}��ܵ�RX�ufGA(���H����5��!�`�x��=��[,���d�ch�"�� ��wY�� �)�/��yM��2��Y���_s+�H:��vؔ]SS�|�8ݙ��e�|i��Eʗ�̛Xl;W�[�����Պ����h+'%'�i�ńi���rVL��%���6�`>{�l���y)���������e�/"I�c�,��G���������l9�A�=a����n�r���{���3�1I�$I=�P�����-H~�ƣ���i03�s����F�-��=)M�z���p���4���(��S����˩����j�4}��"q�_Ces�����PD�����gdC4�۝צ��D�%�+�G����/�3��E�
T5��<c�?�����P_&�Y�	����M�F���
z�������Ӹv���I��� ����2t�c���>k�\Nh��1)�CW���r������ 	=7� z8�������~p�����WB�Ys�۬��,2.�>��$TA�xB���������[�$#GGG}�"m�D�h�LEŚ��*��1_�E���[Rc���3�c���_�6}n0}0d'AT�(�WSCѮ�0�p�q�48����nb�NN����ʆVV����z�S4S��?�{�R� �斏 �L�å����k��==� �x��z������q�a��r/Z�Oƪ�����lm��m��tt<��2q'��O��8	m�`b�F���{���K{Q�A2�{(S=���
�m/a�&43o����o9��N��]��#��w'2�P!�[.�c���mȗN�"���߿���!\�k������r{�����+��T�q�݁�I� �n2��>3���|�����g�lo��>V,}x�T�\���|�\��5#c��&&�q�	n�x��JFC
����D�������|�]�z��(,,���dΧ�!�u��\^�o�Xm�1�a��s�@FiǍSa�"�Pm�R�[̖KA��uuu]�ip�=�f	�MD� z����r�M�<|������q;.쯨�XklkLʄQ��/,���ǭB��벂>�����V�<����/ ���Yۖ��Ⱦ�K>}+¦��"̴sq�*��}K3�%S'���͛i߶μ���"/uX'tL���C�O��_0�J�xF M�ͤ�a�ޡ���̶���ãy��B{;::�ʴt��&㫉�U��]�]��K��3�w��}��]�L�R�ڧ"�����4y���C�@����1d;���x<��P��h�b}��9��A����5Q�5Qg��$���099��ߥ��]7�a�{�X�8(v��޻�;�F���]�J��ܨ�r,��*�Z������������{��Ԅ�#ɿ7��Xa�y�%� �q\9䟖	D�����s-�͛.�i�v�E��o3��R�~:�}�==T�ɓ'�W�+��s��x�Q�V�lʜF5���O�3��<��
���N��&�BuM��[h����?ۋ^���+6uw�V������p���@%��?�'5ȫr%d�i+��/##�a�d�ˆ�N0B)�����5��!�P�{Z}�ZC�]N���H��y&+��~�	��?~D�rr[�{�N�rj �����Zc�������d���� L#���(��m~�/久pg��[��NCR�����Y��B���)�o�t�v�1��)����6��+%�2�!�Z&���(\SU}��*�h���";��V���������t?� ���� p�Z���.^?���"��fzv�ET'LL�˹��:q����,����w��}��޷��<K�ΤjNhy�gh�]&���iD���FT:���e//��(�#lx�e����������񱱵?��Cq�;V�=~���H�p8�	�Tf�C����'l��rܗ�@&j�Ͼ(7�nĉ?��P*q�`��#dP$095u9�I��;}�G3{��Q{��y�m`H�KdH�`��>�W�xC�����s(�ٗ'l�
(G2c���\��Y7uw�c����RG��a�&��b��fP��+y�	���="22����M����X�{�M��8���B��{FG�|�}�P�zWw�0��r�7j{��J8�Vl{����HK��qqA��ښ�A�q3��0ZXXd|�r ),x��#�_
����b�R(r�l(I ���<���(����Z(��ʍ�Ok��ځr�]=�v�������υ�m��~��"`@b���{���Ǌ�����O��dFEEEFEU�/������C����X����I���K����L�����3*w�g��~dh�%K���J�:9���� �n�'���ė�z�BS1�	-F�wn}<هF�o�J�w������y�D3��{����?�9
_���vO��[Yc����3i/�kjT�QB�'8"�ۛ�"_�:�o�݁��$���&T�YH��/X�"���}o'3����a��
��`9CN�Tӝ��+�����_�����z����;d Rhi) $`��%�����˂���[�w�+����V��sUm����4��aی��W9kr}c��^M9�:����D�L�w�dn%j��AB,��BR ?�q���|4C~�6Z�0��̀�"^�f����Bo���`*jhn~
t!z��������U( ����O:םo�&5�q��v[�P�,��k� '�żc�4������Cn��ܫ���#��Jѷ��� i�g³��ӕ�Ӄ~*n�ɑId�S�\�ʽ����$W��_��zyOETC�ж'@)Fp�r�I�99���n{ �h�Gf��Utm���C�ܢ,��>��q�o�w���/��綳)픟68��n��Lv>�,8x09�@%0��TM~�*�"4�����k�w����-=*O��d���b��+�L�7�����ݖ&G���}�I��H�Z����9��Z�=�hoh�����=�~r\�?�C�1}�
�w����X���44,���;�1[�	�C�|n	�H0䒪�j��5�D����Ba*�[�[&H����.�;w�P��j����菪QDN�t���' ��އ�
`�U>~����O=:9Ay �����ւ����ԌJa�m����F�X�*������udW	��
V�{���kjk/��չ������΂ܱn'vY��MEDaڂ#�a #߾}QEd�,m�Un=�|�pm��f���;�#�^olieU������e`���>��"𳧻Q4P3eQeazo:��Lŧ��Q�Uh!�����_�J���ijialIu���f5�X��6[	�}�1�m�6.(��&0Y<��8��v(�
�-����H�G�vvgP���N��tg��l*��clsI冨��v�.�ѯ���.K4�622�
����e�c��!//��g�anO���j7277�Wx�� ��_���ѣӌ���&�P&�Q�8����X��l:4t`R�4ac���b��̤��;�������V�l���������W�T�Ԇev㺡)�G=vVV8m�L�9��F�xy���ϰM�u��RXϵ��so�dl4��M�W�>�s$#�0^���I<5�q�z���_��Y)���̶��m7g73ڐ����9[�ƙc�Gp<���_�����xH�p\�'�
q��7~�JH)7!��^E�f�C�����Z_c�5���A&Ofֿ�!v2�yV�DCp�)�?O�~ѵ2�0�2�K���'G�^���2A?U	��b�A��qT	�	����ge�C�-�<���h�,�	  ..��Ǆֻ�q3�a�C7jdi�++ܣ�q�<�_Q����3��,�������L�e��l�P��i�z����8_D�#���Zc�YWk�8�:\P�F�!p�	��#%n�)ɇp����uu�0C`�FΌ2o;Վ�N����|k�>��jZ �B-0(㔣�H"�\dɱ}
�rc��(����	D@��n�N�\7���ŉh��@��r_���;oУU��Vwǔ��${D7�7�	H+�RKOuUJ����CΓ����R@�|q:�<Ɨ���ٖb�9�7�g���QZ~@)��L��;��X�u�`�v@睝�'��A����������mmo��E���p�b���:�+cI���,���f�\p�T̌~v~���J	b�Y?���6�� ��T��Q�6�k��[#�h��7���wy�
F ���@��t`�s<�]!�P�@1���]�.p�6��;��͗܎S�D�r�ރ����h�H'~������������u������A��+��E�y������v�*���@{�e�����LS�裞`��Lu55�D�*7F\����"=���]C����ԗ�����]|9�%�?���7*��ª�½D"A��ރN�Q�H݆z
3�O��,�Dp݁c�\���+��U�(���P�g��1ۤePƯ��	�{�bi6�N�(,H>��J��f+?�H}��!�9�p�=Ϗ���j$�l�2�_�f����:P7��\�܆4������B�����d�1סe �:LhaoMo$/�P����>�������$��u?�!�zp���p;�H�%�6
�T\Iu"��皙jizm��Tn�j�[qb���j{�V�.b#������~�-w�s�j��
������w�9�#�E�]@˵ƍ�;���s�T�R?t�c��Z=(��]L��{����@HPS�?�xa�n%� X�ݖ�;s65��&&&f熪�ra+7R�3lM�v�E��;�(ή���%5�>sƑ�+**��[|��
��pjh�1۪���� ZgQ�ƾ����rp��3��x6K����f����x�	K�� S�1`���-�Tէ}ɯ؏SP@�m���l8������^иQ�-�"���R�$QD��2XnUO/��USZ�Oȸ.������#����E�(��[�`ڨ�P>��>-F�Ipxd$��*x?n�����Y�ZS�[��$/�y�w<k�+ww��a�?xQ ��(�_�L�w�^��}@���{	�mjjB"��<����Y�ڪ��>i��`�-���s7��:4#v��Q�#.O����ʈ��1O��#�R�b���$�痢����k��o�b�$P�m� �o����`)5�̈������_rs��Yw/�?��"�T�sM���x'����������Ւj"x�_��4Μυ�X�O���v�e�4���:8�C�A`�l��F�쁔��trk�����Dzz���0�z�E��/�.��rC�"	z�=������ &T�y;��_��P���:�����e\�����,N��n���SpEK�8Y���$�����.���3s+����K��"48_]3؋?~|Fj�Q	f_\��$�B�D��;ղ���<�YK?��aF��Q��&�=�j�bI�t/��;(À�'���տJ,�V���
y�A�s����������N���0�\=JS|(wը��s9r�F�'Tt���6��gDΟgDN(\(�:Ѝ4���ލ}/�箢"���ڀ��V
g#P���9E}�>�=�s�����>�b_i����ϯ`8���/��ˌ���`�)�w!�j���إS
��1�UL�#Kf��nt���e@CL�0;�F�)W�E9)TC����}���Cc-8��ڋ���tJŪ���(��;7��ӛ����'�<T�Y�Բ��&���*�xΈ��
�1������A�fR]�{�� ,lܳ�wu249f��.�[p�vе��$�ɬ�k��n��)p]ktZ���m�!����h]��YI��ט}s��,�2�8�7�Y��MKR�R�]�n�r��V�Hs�@��=�H3E�h.��L��><�f���[\�|�-A �y��,���q/�sf$��~�Mξ>M���P2�'М�����������y�b��C�[��^]��w�K��s�$�_��2Ϗ�ͬomp�.�z���2��3�겓��k���=�����A,m��~-���W�Fxp�J-h+�1�����I)hA�赁�X���<�F��x��ɓ�it�i��s�x��l�?H��(�U���̝��+��������8��tv
�l)���X��}�_tr�7O�qq�ؖ����A��4��8���q��o����׾�#�s��k6�L�=�f���	��x���h,;]hG�Z��eu�Pey S�fJ���$�%?�Z�b���1���2����~��Pn��t��Uk�@J���X:Nž��/��Jk-�]��~̬�՞k��a���o���=^`�-M�`DC�h���*�G�ҽ�'Fߢ�w���K%�Ŷ��Gvj!�O�ǣ��S
��m�0�`�@�	�}�Ik�ϗ��)EK���n�e��^܌.�!�
0� ��d�$��/��<����#��#�JI���������D�.0vh}�9#��I\o�AD�ꦒ'�YS�@�7��gQ_� ��.@�~D=n?�������J�~��x�,G5
���A~	��H�U
L�ag��!m��"q�,�+fh��	�9��A6�ve��ϟ?+�?�^[D�Q�����2�8�t�_+M�P?������m�2�j�E�G@e�:�#�e��h��y�l�,"r���S�0�M}��3b�")�D�Y��S�Fk�h�պ��IB���U@?�o?�.�5�m�k�+�P?���k��lђV����m�/ZΠ�w&m9��f�o2Ƕ�ű��/�E���D�w�Z�R�ȪS��z>�|t�.��6ې���C�|�)��5Qg�Rff&�@##ٻ���U�{s&4� 0�(�1��r(N΋#::}�5��O���C��ѡMkd�����Hٔa����CD�oHP�K��H����ƊVJ:����]�	BNS|V+�����k&12n瑯��AB5��@Ã~����z�n����z�qf�rvى�L���"���y[��rdll t"��7� ��6c��323C��G/3��8��{�~�֕�Z���J	~����9��O3�S���Ͽ��m��X�m7ڃ��X�G�̱R�G��v\�\>C�@#P^^>JZŠ$��k��\�Xa�)}�T�58ྈf�d+떖���\��f�V��$@l�KW���G��hI>|#�֟�
 �8��=VD�Bۍ�a�g͔�^�1��(�m����/�oa�m�m��l����yQr�	�t�6�~?�n$:��&^��O�}�	l�����:Ց���%XJ3^A���30,�iR��	fv�Zܽס!�((`��P�)��>�����$�^k�h5�b�C�����!`����mv�8z��TP2�C��8R ^W>��e3��*T��4�鯖��魅����S����)K��(�^��P�L���Fd���Y���[���Ds��L/���.M���a� �񒠽++t#�N1�%��>Y�d�V��@�T��eV��p7��nʦ���O�_���k[��� &�~9ʀ\?�*�W�(I'���H�~�/�����A��.��xl�bѫ}�6�^��9��h����u%�a8ۺ'h}��kVؘ�s�E%����A3e3J� Yt�ћ�E܀�z�1U�V��8e_"�`@��� �K	��_%Q5rU�^��	}+Rq��y�@(�-:'��bdY���R�fZC$�F�̃�WzS����� ;$��J���*��Fo���ۊ�fMD���P��OaO4tqȺ3C�QtF>���m?����� )��2�
T��n�%X�R�@�3�8�Z�hY���.�ʹ9;�B�Pq�7�3��9�w������U�^wcT_0bs�l7���PY�o�ƚ��:,��I�(��D����K����Ef���O��{"V���gB���l�؋$z��A�О$t�E���f���*o�( *��&��I�7&r(���8�����J��`���������4|9��?%׉�+�~*P��9;X�6�ѭ�pi#ss�Q셠k����#2�};t�Q(z4!��J7#�@_�/���Ӵ��p�?
�.�����u6JNk������ �y�	���ի�ɽ/aw��G�"�{<Y���1a���WL�G{��+vgZe�������*�o�3|���k/�3�h��&A�2D�Ñ�l[�����$��WE����Awp˸B�[�<˅v��­,����<Q@�.$�p�6�IB����"���0|��,8w&4	<��<£��0���K��X��c���B�Q]�sz������q@#��L;�� N�T��1T�pc���h&���0�$��lZYg�ޭ���0@���`T������+�X���D�}`n�����/(7ZD}<���nT��X��vF�$��&?~,O}�7����7�T�d���ޗN]k����k˓����ԫI@J�� ���@�1���	� t�
y ��cok�o�4Q���G3�7ʺ��ܤ��V���w%�i9�'��QF����KCW���Ǉa�d��D۔!�w�7��wJ�/<�^щ�ζd����E�m,�6
��7F=7髦��b���@܅**1�R�Ƹ��e�����c��J��@UC�R&~�rS���n��]Y&l_�C��]Bve4�� �#o �`>�l��š��03c3�&��MD/�244�ZQޗ�����
�I�Q����-~�,Z�C>4������]��BVt���uh�04h�r�N���N�S����!��?@C��+�;�����+r��J��\؎�J&���B:��h0�`Nǣ�����9�M�DΝ;�%�W�,�2�%��X�wb1����<қ���`T)`�]]u0D^���A������$�[���f,��(O��J*ڃޔ�;��ʊ��� �Q�p�n��ܠ2��`x0�)�)r�,r.�&�nA� ��ab+m�.vL��;�h�sZZ�NN�-iwΚ��B/É����5��U�q�jx1J _FGb��т	�e�㑿�7�~�߈c��E,��;���}�N	PTTT��Z�_t�Ooj��^2֙<sF�5�e�L�L2��ENs;��pw�����ԣ(��--��{�7�q`"E�W�Y�r��!�;	�(*��r���HW����זa���0VD9γ��@���ѱN�����]�P�c���[��W�-`^�?A��g']���<r>�𨪺�^,���`��uP��A(�+7?�È����0��ê��q!�F���p-iU��̒g���A�y��`WQK��)�� -�|��~]\�c>;"Yp�l8ۙOh��;(�<"��Zo�8L^4��������De� #���Zl�6~@�� �hϣ������vN�J ���3�����4�a�xs��D��(�`��g�~ʭ�*	%,V���y�&��<T`�ѮP||0R�T� ԇb�x�=HII�mH�������*�u ��Elha�th��sPST�P���E���8:u�E��Y��aT�F]H=��^o� ��ާ��;?���N�y_JkAC[ h�?��gKvr�u��0��c
<��؟?fAܘz}(h�8Zio�2��)`.А��;g� T���H͡eD+ШD�齂N\�0@�"� �E�:��U)�.H3R���D�����56�\P��g6&�����V?�ۢ�w�@⌌�C��P ÇH�-�8�Ld�R�6F4S�?��ox����p�����f�kc����������C�2)�@=r�+�y��䵏�S��r׊o�4�����wc�Eߟ�*�v� ����՛�eM}}O����'[�Y/�0�������&s����E/Ʊ��VF˷`��������y&/�E�UX�NLL��S�ȿuj=>�w���Y~�Yu�K��f�q���\[_���EA����݅JU�NE^qN-i�Ҋ����Ȳ:���H�6�'j��RYzb7w��cL������宋�.l����ω��dZ��c�U����ʻ������wf�����!��n�[I^9M�w?}��t��^_��5����z�Ћ8H����f�ݻGxV�YV������..���iسaǰӭ��챇_o8�x����b�O��ʵި$>}l������)�%�߰I9���fǤ�{�=��r�(�X��M..N���^����)�RA�;v�8?8�/���߷�ޢs�oA)�}���)�,����.\u�+��pt\�Q�����l��_�Uq�'"�ٓ���)�"�(�7�'�/�Vl�֍�����
febd����ڊ\��7�p���#�z�W�n�J�[j�0Xɭ��&�fc]��j�pqƆ����!�{KKK���d�|�2s�P_���΋s���055}(�޷�G.lp���ؽX�4�䩃��500��f��N�>��ꡎ��5��_�]f���~mT�8|p~�Zr��C�������o�/�b{0�I��>G�k�0-g7�#:+���U�D�J��!����GF}�ju��ċ��u���v�����kF����n�Q�_2�\��&����␫�i��:9������MHI��Z�r��0p�j_��Ծ+v76;���{���Ij��g��W�����$O���5��
ꩬ�W� ��u�
P/�]�
�c���"�������o~k��K��n�-�$����o���D����t����Ф���&�,��a:xa��ę��%O~�'�`ns�~��~X�aF���	*p�Jb��nLn���SV������&:Y-�A��A�z��m������ݝ;wVF���i_���Ż�/wn��'�:��7��')o{��R�Ͱ�:�ô��e�]ң
7�|9)�z��8ne}.A��؅�&�<;�X_��vd�j��~Z�X��ߺ7�w{��������~���#R� �T��E��/�`����X����T0��C��{�����϶Q�7�Z����	���|b�TZ��O�f+�!��Ɨ�eb!�?�/N��xZ蹯����4��컰ї�������

M�#�,�D��Vo\7�\6���Zy)��m#�M{����ڇ.{���;�Su9��u�7�N����������[3���&>�LX�v[Cߏ�z^��S\l�SU0b����`�l�'�͐/H�	yԣ�,..�N��b���gJ�9Q�qA�֒�t�J����=A���o�]�{P���;�(��xM�ל�����QgM��>���5�?񝸀���##1L���v�Pr$v�+l���a�R,��4��-�������S����7�U�$]�9{��go�c�j*u��n�؋�<1����K�����P*�9��H�ߏG��j1�/@ڜN(��8�q@�@~R�W����������r��^S���P������?1�
��&��2X�8۽��vo�ݔ�l�F����ʇ.�T��s�e������k���7�����-
�F\s��֟�Cپo��3���^KHM�R�(�e�P	�$eˮ�죒�V������I�b,%$k	S��l��3���������yK����<��~�y�w����ҫ,�_s����^_�4�G���#徱�O��'ﲾ�K�!Mx�"��߷�D7En����o�ѐ�*�1P���@�*Qݎ��"��Y�D�X-M/�t� =�ssPY����\��������XO���_r�N���T��,�iv�<�P{.j��CO�����0�����6�y����6������a%��TMi����n�+��!Bp�ul`e[���Gn#�ߐ�_	tq|/�0/��6�yA@���?t����k�v,�� �쭭�t�{c��A'h���+�����b7�w*x74<�M��7&��dR���)����%Z�d���Ϙ	��P�+��}RM	�G~TVv�먮�Aݎ��K"�J��UG
ۏ`s#�6Ľ���;�=��_Hޟ�`f��|K�������2��bB���hpc2�19�HA@@@��� �K���L�K���c�	q�}��P��W*��9`�Rw�Pn
��������^X��꿳�[��UZ�#�3��"=�~ȧv��A﫡�oߊ-S<������~Wv�-�<��G*I?��n:$'���lUSs�O"��۳����1|Ev�O���mZ:�,�1��C�&z8�Ŗ��'���7����'b����(Q��7,g��+x̳t�]��`pc�U������{S���ް6M,'�/,dx3�P�sb�N���"вRP��`�]7���m�[�e��LhL�(��WN�	���1����+߼=�]��JVH�V�Y7'�����_}kpC�7����6rk�	��1ֻ����'�	�+\C�>\����L�	j��DM�s�����
��a�꟔�4���8Fs1A"�ߒRx�R!�_�~X.7<��iV����(Xyw�@�t:�R����r�M�����Muԏ�J~Ք΃����ׄİvC���t9v����Qq?�_��
ݒ�9TGp�tl����oB�X?��'+=�����(���^�>�����aF����+\���ka��b�;�o����֖�"�ʎ�X��{]T��^�'_Pn�7���/xa��r�]��%Z�iiK�;n�	p��mݺ��0~➭ U�'0L}{��y�,�İ��������U�|�cN������xZ�Y%A\��e��&�:f�#�`�|�ɯ`3=�Buը���?�GJ�U��xA�u+���J��@M���V�������T���U��!]�����Smh�`x%,��K�}���|�R�V�v�nk���yp��U"���n��肕�g�AJe�l�����*��}o��g�����Ư��g���Tr��'�A�.�'�5Q�9�[v��ښ���O�=�����=�v�y2�7�]R�sq�L7�1�J<�,���$WK���������Pm��9��1ڦ�^�9F&�����:�j�!�J����m�;����Q���+vVK�<�Z�p?Vf�������t��.��i�5dd��s�-��Haͺzz�BBBv�H[S��K嬕�nf,��_���{)BdGGG��ؘ_A���D�_y\~���s��cK���T��X&DvZnL	t#vq�|��dhXX.Wx$���3��������t?��������1ע�����l����8Ḱ������)��8�s����j�5���
�Z�3	A�ao�#�K��QCb �(�k�94E���X�7��-]�Q�+��բ�JQ�~�ѓ�H�׭t�6bC�s.���c���Գ���-�(-���J6����d��1#X2&8z����.ثn�Å�d=�>h��&��zN_M|�����P^̡���")n�����2�x�pՄ�!�ګۆ󩪩҉.��3����7��F���(�y)�͘1t\�c�I���S�|�qq<q		�Z�BZ��ҽ׭�/��G���i�v���	7К�0e%%_Q׃/B���>�l���=p��jFUD�݌�Us�|��+�����_:�I���X�M�^�\:����	���ַ�]���#��`(�֐�r���{�/�e���T�k�ช>ܸ�K	|.���۾�^�KD\��m���=A��)���������7ov�֏�L���?�aR�!��\���h��R���Z[���D��ڠ�4r�=��m ��אj��xUY�O��![76����B�p�෗�gf�ǓVl������8��e�ܞ����X���:\ʙc��
�+w�|�{x,5��9�J�
���֞@yH1ݣ��x��A'.�Wܷ7�j��� ����d�����5e@��^��~��@\����[&�]�x��4�V˯�9�!2Yvq�����v�Ct;��`�&�m���H-�������W+���988���/�k�ψJ{�.T��6\����K$��i�m����#mgl�5#+���<��iR���c`��)\Q��M�~�2r����s�߿;��߉�8ߩ�e[b�Sʂ�6P{���Gy��a�Nrck�ث�i���	�۶@�K����u�D�T�d�c�� /�d����?��4W9�3�F��
o��~�{\���N$��p<%Ҡs����9UGUl���[`�oC�	�^�x����x�ӃƻKI�KI��k�t@�F��
����>���?�F��u;�D5��fS'��"�G��Q�=M>q�zFi[&i̤��wG���w7���RO�T�*�P_��-�-R�|�d J8G;�y�P�ap�}��;�e�Fz��J����H44��=U������ �`'� !]��t�:V�-��Pd�j0�]���tc�2)�Mc����t��(����x�P���@��>��vF2?�0�z�G:}si$&�3�z{x���J�h��	 Ѐ)�Y�߷)���}�
)�NwM�UPZ�R�i-_����~	�dm�VGQk�C�waW�������B~K�uV�=��Z�Ýy��a�sn	8��-��v��(�?fV9d�4�K��wn��	��џ�yk���_��76�Ⱒ:�A�3���ONr��Z
|L��a��`���>�c����jMąƻ�b��+t�U�0=w��yߍ�4�)�n���v(�M���/C��{��#A����W���`Ej�"tZ�f��2�����.����>\P��܏�[�s6x���2_��ͥ/y?}C$Y�3�]M�R�ƙ�����b]�x[���98����`r�*g'{I1�xÆ��!#���G*cETj�H�s�X��^{�ޭou��x�3�dd��:F���Evm��4����������*k��X_>t)��ASW������k��~����\ffe��\�>mOCM���-hZ���B��j�����#��4��RW�03S�q�F�<zT����@�L` �}o�_ j�:�k˂��SIn�g$�>��^�BK_����jU;!/s0���wL��.Qʱ#�o�m�h�#�p���S�������Ƽs�_�ͳKs���xl�V�Q���...��o�#��6%��6��J'lg$��h��v�ŊnN14y�n���v\����K~�l���w
}��衵����߬�Ԑ�ƾ̜�^������b�J���M#T*��GGVƇ���橷pv)���(��3Қ��ٵR�t��R��/�u˺���ݽM�c����jj�em��ܹsQ;cG��^f�մ�܇�p����Co���(�29�4���vٱ�����#��n�LJ�s4�)�z�^�����U�Y���x�h���ԙ��޳Z��Կ?��`��p}������si�Ƒ��/A%����IkO~�-�<�B��j�:�LP�Œu܅	�C(���ޝ�!��.V�u8��٭d��7��s���Բ��4��J���vN��۷�޲���G����~Õ�D�~м�����=�?#�@\RRty��VG׃<�ssL�Ca��l���A{�_C�z+B�D���o���/'Q���wr��ּ*�{>.99fi)+לB��>  ���j���ȍuY��Q��`4K��\�/`d-a�Obbz��J�O*�1Q�Ū/0�l������x�����8�w֙���U~�T���*۫�X[+�{�g�����A*CBC�76�w����܀]�yt�r*BͶ8����{�2��T� ��ɴ���H���@����h�3�eJ�1�]ȡP�g��DRɩ�((-C/�E���%=�Y0a�{E�5;��x�Φj��3Ԯ�H��V�ٝ�F��F�qҰN�����?,�*p7������Z�^�&�sPc'�F�+��p��>'$�$g>���"\��Y���ݴ�������~Y�з8�ˠ-��^ύ���c,}}M�����<;@��~����+���q,e��<ڟ����� ]^+`z�Z�ԅ���g�G�i�<�$B �����\J�U
*7�Kt�d�I�t5�Y���g����]7OWݽ�(z#���4z�`�qQ˷|ٽ���|�Wq7"c��+grJ�l�G�X���T������<�+W���~?m�'�5z���� �#��\�y����w��R�c�V�桡��#��H�O�����S��bu��a"��ח��n�����W�2z^Hf��r�T��!Wt�7���$;�tQ@\�sQ˃���7d���^�@H�H��	#M������'S���e��ގ�_�F��섴v���[[ge�u�0�
��R`��&߼�5Y��_��:a������h�����O�V���R��j,�c4+��1`?>e_����1��ZӪ����9�������Z}0�؎��w�gG�X[[[zxȻT܏���n�Q��/BOWW�a�pCR_-	�������,s�[���P���qQ�#��3mh�W������o�3QSK����+� C_kK�]����s9��8p�Xe�F��hmu�-�܌8���/X��'Puzpy�B�e}�̤s�Y4���6,)W��MP����w}`	@okk����O �������<R>�uvI1r���M/��=8LʎꢧR�h��{	(ϰ*/�n#H�T�Ԏ;�x�����w�DE�ntȿ�LW�<ӫٶ�.�h��Н��_=��B��4���2��V#��՞n�;؞�1���T5B�\
m��Q�ɓ'���=}~V��t�5	�#��]��v')Ů��٤F,�trc%�%ҭ�~\1�tv>ەsY(==�▼^Bj����Uo�؇��?�6�A���"�5�H�Lb��)���:S@ڭR!7f*��h�2}t���y��'ǰ��V,��L�=#�t�� ���-=��4�F}�zn�ϳgϓ���ΏD?Y��(�N!ėC�(!��J���mo�U!��q�T�X�4Ə���Ug8Q�~���M;���� }�K��4��z�Y���ѩ�sD�H�B�����oD1���@�v��KyVS����hv�p��[�e��Nj6���j-��
(2�7d�r,yr�=��B���hԆ>�4풲��8��ړ`��.����.z O��n#��̬/�~�u�N���U�#3Mht����(H z�:0X ���B��-�^�$+ۮ��G���'~Ɉ�������L*�Gt�nI��P`O\0E��ys��}�k!!!��폷n�zJ)9�$��&M�����8�A��!�Gk[���п&��wo�[9w��~�]�y�MΡ[��=f�e���G�����G���_A���Uz&S��塊��z����S3��=\>��-T�s���G�o?�E�=}�4��bc1ף��h[�3��u6I�{��g���d��݇j��x��b�����o����츢�@�_u	������Y��e�(e/*IJ�Ex��CukgD|���0M���%:͉�]c,�#��mU(��gcc+x�R%��ԄGk�|nW��@`n�e�OԨ����ц����V��P���EF^;qQ@���d����lg|�`�#�sO�q��ot;�����b�O�޼����|�5UnM;>�qF�u{Jҟ���I��ƻ���/a�l������Av���hЙ��/G��D,�7)�rA?�@���1z�u_8Q����|�X�ڲ�a�)P��	Եn��5]��Ft��
��b ��HL3#+����#�^��	���c��Z�ǸD��%��_a?�m"�]�h͇VQOR�`��k�3�P�e�*]ũ�$�F�7
D����
ko]������Db�q��LM���F��H'�3S��1> G�9|���&��+��Y�?��_~���l�2z�Y��
���r|&h<����Ay!9��2��ʋ���#����
��ht���Lg�s�V�^�*:�bE�C�j��L DD�c_���,��s���9ϑ�0�ø��oi��G��4qDZ��I�gS7w���[ܾ�z�<q+;{.�Pۓ�a9�r��r����.J�,{���i�Њ@�B��	`�t��Fx��� ��Bd_��<wpV�c���N �O��;�t���D5��uv#S�6��(ѹv���|1L	�={d�z�0(���k�sjK�lq<;�>�D��j��A/d�  RE������D�x�6����ں�?���H��_��ǞB��܄0�(��ȁ���t�ltt� ��v\6^$Z[_x�`r[��_�����ėdyL�=o#� ��Qv��u���7�ޯ�����|(�X�ȉ)Y�&����_1�D��Ց%����'�y$V�5.1ѕPp̕}�d��("����y�)P<||&b5\[:���c̗���1��o�#�-��l^)�xxĉL�d��"N���R&��^���]��[}؎t�X��G��Է�`����H=e��n�/<�ָA�rRQZ��脠�F��� ���GC~�M�ڎ���`j��n��?�E �	��4>���_x�sB���?L��g�\O>7P�/*�
:�K���sn���0�Hol��*a�Nz���0�����	j����W��0��0}��
�rQd�j�P��� 3����V�]�QCm���m�����5�y� �����dp�
�)�ϟ?X�am���Tԁ�xb|����Ik�c��r�-t�t���R��ظm`��%�����C�)F�/������pF�_��� 7�㓩/=��~G4��4k	�Ig}%|t�X6�~�%A�=�;�s�����`�-/&	`�/���-ii����-n޺U���nc*d��uz�8w��kQ^�1uN.�Գu���-�p���d�77_�uo�tء�$H�L��Ҩ�y���3>������ƺ��P�騮j��Ww)S���X�p�o���p��E�P{{����i���C��*��=�SomⰮ�p S��=
��cZ�Mۇ�ŕ���0Py��p���-�|(<Ai�t�f�o����ur.�Ǹ��ݦw%�{$��K��ۮ������<��61{c�>'����oTTL����������b�w�&Q�i�h����/h�R�դM�s6��O���좗&���?O9-_i�by�@��4�H<�Ua���U������X����>��t&�g��6@��D�ĥu��,�c�J��9�K��]1���j��?�E��![}�[I�(��7�}J�m�w��P�����X�9y����S$�>���G�ߡ�A~[�"�)l��7l-k�u��� ��P��w�U������pp�Er��[�. �����\\\m+��Bt��F�ز>�����G^_���OV�_�������0x�@�?�Z�֧ǭ�r�Ŋ�i�tvI5��s݊�T�%0p����vyujzm�-B����L�ׂ�j �er����#@x��~��.j�@(��^���������g���vg��w�WM�A�}#����v/e3+�1�Z����wR*��
7ޖ��zz�@�x�nG��Ok'k�lA-B����M��>q������VC�����~B��L
7=~Պ(}��J�*�!1Ҋ�X\Ӣb������bX@��2~u}y�8�|�{ѹV�u���J����XG*��k��Fj�ZaT�������mċ�_�n!��/��%��zH��k�A�1fbh8N��=<��b�^��_
[ppp�yCX���\a&�(���׽�����$v���߮��k�+~�V���K��Y����XZA� �?`���Z�5�s�������wɊ����]��������{�õ��Q5>3}`�.%W��x�!���ah��ŧ��\T{�*�}���$�%^�0љ��K�2pŐ��<3N,��O�c�s��'�g���S-TN��肬�ᕠ�w4��� |���M,O����)�Gl�*ޮWbR��m��Q'���0����W6���^g��P�A�ر�sjk������Q_��Ovt?�ʣ���O��F����q[5��V�5wC�!��%��Zj��ړ��n��a�0����"��	ﾲ�2�z!<.V��qQ큚��yi^Ŋ���Q~5n<`�0h�����L
e���-u�����s[Cö�C�g]���(��"'�nˍj�i8oed�$m8f�j�K��@��>�Vy^��qdE���8>� A�@X��In�`W�ĉ�9��ų��A������.#A#p�}۶o�90�_��Ý��({F�0�9�R�t�'~Gw�W��C6�����AIi �yD��]���"�.�̶I�K	���[�������l��݃�XV�Rv+��&^M��3K|�p�V`���t�����8��h"�~b_PF�o�k׾ж�ܰ*�$�`�{�+D]YRv�K;��n���2�	�����(A�A+noG�pОm�L���G1�c������6颫$7R
w�������Z��=��2�"E���bԉ�73H��wڞ�G�@?f�=�yAs��?n�k�!�>���h�ހ�X�8����max��kr]ϲH��B;��%wG����l�&4�������%��}i��=�A�+�4QDih��-�1Xf�0��~0æ��)lR��;~�x�F,'H;���y���X1Z��ʅ9Wd������m����ce��un�^��i3�c��>�&��E��{��°����b�3N�<}������1>�k�Z`��\�]�^:[ƾ��%J=��ú�R�N2��}ى `t5�"�l�n z�Oa�xm"i�M>zs�c�	�:�1��C�)�o!�.�[�p*Wg�L�L����rs��~3HZ��my���]->>=���0{
ɋ�����<YɸP�'�}@^����U�jC^�y�r��P �����wf5��9߇+
�K,� �K�l[5�)?M�PĻ�٥��+��y���	lа9����2��9��F8���SfT��aO�o��0����M��"��E7�&R�+� �s��ǹ�1�Te�wnt�Ӈ�HF#��o�;�Hq
`�R���|����̉�s]&��g��T�t�j-�2����d�I����:R8L'zJS�B��q�#^e/���DgN}:�R%I�:�۟�{��c��?
I'�ʦ�3o3&��o1�o�u��sͼ���2��m��t�s/az+������}͹� �ii衙ϼ�e����/�*�x�:8Z˯nNB��U>dd��j��՟G�ج��n�x$%�K�&~6kg���_� �uݏ�����lEP�7�\��N� 4�ҙA�"
	���6�3q\w�m�=!�qκ4L��f�ƚ�s�W�a�h�@��T���f��v�4��n)�;ww���YI��)�|�����ҭ�֛_ �Oc�Q]�n&3�տU>+,��3n�	ޡ��B�k���T1Y�	�W�pG睵j�� ޥ�9}�Ѽ<<q� ��{��W���8`�An���@v�6�\��i�c�z'�.J[��fX��	H�A|o��Z��y��s�eԋU}��E%>��DbU���D����[�#H!�S5;�>���|���c�`��Ũ���D6�1s+����Wȭ� ����E��q�:��r�u{�^\Q�HgMy����󝬰�v�.$Ӟ��"x���%57����g6˝�<���Xa�*
7:�qfo�7�%�?o<,�����zf���I��},������^vY9V��	�(|ͭ��"JPE|�!Ӏyl�2���gC�S��]��T�n �����R��Q��S��nHd.Wx7�gʴ����릔�����!K�u�T���i�ܯ�X9L�@v"��V��K5,mЌQ"��1�x&�%s����wJ�n$(�
/TUn��PhGv�Q��OwD��?���#2д�h-Ɗ��t	�a�N�����_�hk��\>�Т	0{����g\��(!>�WD���@a�j�֕����c=e0Pb���3n���a��7���D��E��Q���|l�J��Ġ��u5���L*~�:�8��~�����3�Q^WO������5�@D~u���yp��Ci�۠Bt���Z��{�0ۆ֧l���Gz�~%����i�� 8H��H�#��~�^|�z����@��J�dk-��k�����)F�M�C�4�}%7��+���L~@�
�w+���$��{�	�~��b-G.hm/@�Y�����;>�k�i��nA,'%-�K(L~���S�j;�4��.���!xf�O��3.����C܈�����K�ԪydV��tݪ]��E��� nT���	6�T�Ǯ���St.x|����k����ۄYr��r���Z�x�O�KK;����Z�=U��!��>o�5��B ����69�&F}i�d0_��VM�pA\?��M�)�xORC�b���:4�dt�A�;�q�(�Lg���G��j�u}���
���5���9%Co�ْ'9fQ=`\��ߑ貕�Bx�4���>V��X�^
����xW� ;$f���'�T�k@:zw�$�����w���n����2��/�QJ��0�`�lШ_��K3�ɕ^�����KS?�L^2Q���:�i/��O�	nz'~��#������g��+�IX+S�`���/��},g�Y�����_a��F�6���]o�T0��c?�L«�z�8��zh��gne���7V��*�遜�M�Q�yc�5�'jo��6�)S<H�fD������_c��4�=�-6l4/^�R�s͍Yr�6�:���T��O���ؕ~E���H�6��N��8g^���T^�յ�z�13}�����1�A�N����p�Z�[���q�w���"6�̮����L^��Κ�<�`A2Ȉ��� �K���d�;drD?�Zz٩r�x^R����B���.']
)�������2��'&��~��Yg]@$��Uwd��n�03n��v􉶓9�W��1�����#Ji�]]]{v�9��W���7O9�L-�̪A�V�EX�\�;�:���_���lgg����MF{�0>o�Kωu�R�h��ұ��;X���СC~��8�:�}5r����s���6�O`fS�N..�W
�cX�5 XrL#�����x��XN���p~�U5g�<#*�W�ֵ�?���Z��].���P��P�������3k-vXQ�:�w0KVFf �i�].U���<�`�9,��}��կ�Æ��oq�,�V��Rҟ̏�Tę�1��{�n�:��y/�7�&^��t�������.��2US��X ���.`�ծ,���+@;1G;i�͑hu�ʂ�PԈ�o͐Gɮ���v���$�M�-��>@���4��@�<P�G?9�yk�)B�^��$�;���{3���[RR����a{{��6j� ��_��6n��5�+�-9N]���&����%O�l��J27��od��ӧ��HZ�r?��	l��m>9s�g���e!�I/�#N�{�m����̺�@X�Dk��7o����a '������=�����Q(	�RD�y�ͺ>Wr3����<jq$9�n����SR"2a�Iz���3�_v-�`'U_��o�ju�K��he']2�^����γVb����N�ioI��&��\�o�:�_Q-K���5�r{aҏ�9�5�v�ơ55��3�Y�V7	���3���ۚ���y�@P����|3��
�ؚ�Ȉ;���i7V�����\ju\���]�r���m��!�9��=�$m���K����ls�f��'b�(Yy~olM"&����E��.YKٚgIJ>�7{��dq�x#/�������}���F#�����m�zc�ן���<���A����|�ԍ�F�k|^�p�om�V��Y��Ɔ>���!L�JNd�u`t4Su3��*���qz�� D��y�j������8l�������{э��0sT�K�D[>`4Z��m�Sئ���K�b�f�L�����K�E�����9N��&�c�s��(�^���2����$g��P�4��H�kV���G�NaI�,����/~+��U}�<��+��µE 1<c���ߝ~A��[p$ٸT�8p0~ZC��ew�V)�FB��o��t�  ^���A�.d�S_��8�Ҝ���-�����vϟV�+Dtl����XI�Z�Q�<��q��҅��ݎ�'��H#�& "}�=�9͎��y����j����@�e��@q[>�b�{Ĳ(�
������6�K����H�?.������M xB��q�ѓ"#1���T})����t\U4srsŻ���u2@��
��v���nf�jr$]*�|��oڹ��o+6JWbo��G��xV�Nk�� n�H�%����5��V�S�MNճ>y�D�)0���ř �{��]\\|M�m�@_;tSV��9�#���|�W��r�Q��^=��^}�2cԔZ�_��MP/}�d�g�넔fh��I�8:�_��3���/9n�Sui�n������F��O���^�*)qD�Y�D������㕌�R26���$g'��H���'�#�~}z~��������e򿈈��JKJ|��u�H�u�~u^���H���6\02��)����T��n�[�!$2�8��겚�k�
�=��7�.[��Ġ�h���h�A�r�e��=�x���I�/B�9��%=�[�wMїsvǍ��z����C�;8W&�@9�Q�ji�������~�(}%��g�k�P2�pƝ�����n�a�5.����ʂ��YD��Z�_��,�@�{1�Y����K~Р�:��Fo��)��':�&�g����)������u%n�_"Z����t�GS�'*�9�0�4o�-��5(��ϋ��Tz�͈��{���J�(�Yj�.�$Ž�_��4�4kd��&0R�pj���1z��Qa�����`,�q)J߻)6v̙���j��H�����&��S�X�T���ߏ��XԄ��[]ȹ?�,�����;����s��C��$5�ǩ{���^K�������/��ء$*#�)-++ہ�K�2�@� ��Q�!7��xV>���-$Q*%�-R5;�C)Y��zbae0
�}�`)��ۯ�
�Ǐ�2��{����r���Lė���X}��oAB	J���9��[�Xc=3�b��\C�<֊lJɪ��DkV���U���-�+F�)����yx����� ��	�KO����,_y�'DPz�B�'�ka�9(9wDaҶ��ާs�`�5����h`��Hp�zK�vy�:z��'�B���_fI��1BH_�~S�s#�A,�����*_-����}ɹVܥذ�}��g�n;����b.�<I�^f;���+�z�CTSH�{S����ߴ(�,������C�3l�M��U0Ӣ8�XU���2��%n�;�ʱ�����  {�"��}]�2c8�o�^�֯"�wu>_<�b��j��7��(�|���4<�ф%a�sw��J�Y�b����Q�&�KjE�Z���j��봜�Ɯ���V��B偘��7����ʮl%V(�<<S�����fF�KVv���V�T�Ұ��[)3#���+-�>[�ib�^Y��&�LI�`x������eRyAA��?y1+}N{)�^��:r8D�[rgg�f�>;�qb@ro���dRZ��yx��ʟUC(��+�̤)Ig�=����ة�k����qXM�8ݎ9��r�d��!�b��}B.t���:�t��{�[��}T/����'���!�q`�eCT��޽{�m�sl����K�<�a=Yǽ�����\&]�f���\�#_�C.�n9�Wb�|��K��@�/P]O%�D]�|��T��+��𜝏�ȻͦT^!&sC��w�:��r&�����L;^+���Q�㏼D�af�(B:�%�4�|�5�W~L��2���~|�<����<L.����Kt�kӨ������@�;�N3�x�a��VG�r�ZWW�aZ�Bl�S��r,?�J�і�� ߝ������W[!�Q���2A�@E����v��C� ���nK����)��+��UA�-Q"�hʟ��i9�j<?��P��r�c~&��)X�>�mb�+y1-�uy�G�2���?�N~'���e	�yG�,i`- (g(����FL�v���ըC-^bFV���C�}�Qa�|�^�!TA37d�i���]�*�;�x��5��Kr>��st�ԫ$N�sIMʴ�Ӭ��u��ϭ�6X�s�u���8�����(�g��c<+��8��9:�z�m�.�kb'm�صp�t���Ȉ�n�D;�׷O�F�=��Zk񲡻�֚*P'+i���Ǘ�+&K����j.:Լ�R��Y��f�Fϔ���F���r|kW����C�(}_tb�n�^��� ��*�V�Xi�u��)��@�q�M��O�m�����P�C?���q�� *�����)�� k�;n��p��!�*���VҐ�FzR=̪��`�2����f��7z����Ml�5�i(�6社�s@G"��W淾�`���ذ/�ᚗ�^"F{�O����P�� 2��tM'�J9Č��vs#0�{�q�<�k��i|?v	��PMO�?�Zp��&�Ss��.�ڗ��j\�a#!�~�ᆫM��Ǡ'{�� `�`��Bj�����>R��$'� 6<z��hW}}}�[$T�ؿ�%���.\�*T����J��]ϗ/���eW��j�E3^���]J�`o|YV�x3�IKK�r�#��֯��3�uW�̖�Z�A�n@$	�IhI{�^�tV�R�y�����ݡk."#�(隽%J�[�l{�އ�\�4^�ٞ�����|�Fn�����$'���0b��ŧn|_��T�
W}׿B���N��7��Llj���Іt�A-VB��}ԠO_J��*�3=���.kU�����[��yՌ;u�p]d4>_�V��5��`O�v� `Cqׂ%toÖG�s:��I��@��
�w��ڧǽ����H'f�����'r�;�;�4J�7e4�)��yR^��?タymn��'���p/��U�2rOU�9냩��J���K�"gZ�WYQ�-�6�W�}|��Į0R ��f̴q&wCR����ѣ7�!��h(}��+����Ul4��{��E? `M압�Q������ڢ�.�������'����i���L~��lx$p� VUl�Q{��P1\͈J�+�pW��o� *i��/ۃ�l�>���.q�X�Z�TF:��^�ȼGe���<w���q���ku'��z���]B��M�ʡ%�\������8�kyz���3�D)`H����6@����23���.cͅ��vX+��i� '�qw�L���!��z�!]s�BS%LO�&�!�a��v�}��̊��ZN�k׾V�׭^��ϣ��M�
��h��9��?�z�ҋ�ڭϭ����nGb���~�d�Jh�0I�rD-�~&X��MoWVF�WFT]G��$�SOSS�s�"L�a����9�G�� h�#v���m,��:���$�!�9/^��?�N��j�Ǡ���]i��'6����q�h8YG?5 _m�¸��>�_YD�s�qh��|�=]Ϩ��!�Y�b!�����{��88L�ϐ`�.k@{d� [�ێ��޽��\p���gDFnC��{�v��$}��KzW�gX@b��<ƒ�އ�싻�����u�:\�H��KƾK��T|:�BN@���:��y�t-�1�\,�����`	Yd+��=ܓn�H�U7��1�����p���<Z�lF5m�^�k�D�̑��Gd4Vi@�F�}_���0skX�5�%?�g+:��DV��'�J� �!��f��Z�r���Nϴq��7���X@�z.C#0�̏��H�����E�r�91I~:�[��?z��x�v��:�
Up�)Y����`r^+Z�w���O�s�7����S�f�N����)�ރ<�)�%#j��h�������AC�ЇҪ\�'ˁ�H���߁��`�O�1��W����C��%N·f��UzP�ǿ@��P�墓�{_��\o�?Wp;hVI�����Hn�/�T/))AG:I1�_�nU�M���B5ڠ�hL(�]'>�'wu��1�A���^�0���u�!o�8��S�ndd�v��	�]�������-5o9�&S.Hvt��u�(��t_:��vh�H�K�9=��۠
W;�����,>9��n~q��jm/R;�&tU��Y{e���Zs߻�Y�yu�q��VUb&�9r�"�h=�k���+A��.W��B.���"p�j}�}�_�i�>�8p��sjI3�.h�o��te>�?/��N'8!�ov�f����ʸc�9u�֞����6�\�[��?�]�Dñwa��ݚ�yϫX�S���e��7op{���w������r��Q���7oޜ&\�mv��Ә?j#�B�_-�{_>'�*"�����������Tty�DI�(�x��ɚ aM񋐌���>��ϸ���\;e�Y�1#�/l�:S�5F;����^X^H$����?3�#���s}�P2:�J*��ζ��6�D��ڳ��&#j�垿W0�Y�����.!�����~ן����v<cd�K[D�)P���v(���c���,����(v�'�Z��
�Y=D��c?��ͺ=b�Β.Գn�	6�{H�BK�Pd�h9� m�5Y4ck!/vp"5�L�Z�p�#	�@�nAГ.󔎟YD�ZIE�����K'|;�#���f:B�wF���z��쬄f� ����B�D���1��zM�vL�6g0��r[�����0���	,%�6�:��+���~�^'����ַ��y�Ol���w�"������V�v3�D����S'�����999���g�mb�z}tb����c%+���"_��%�e����-�yé-�\A���j
~y@BV<+e?K�:�>��]16�݋_މ��ҏ���UX��m�iZ@[��`���%���%%�GC�A��N�j����]<�[�L�.��~�׀P:��F�x_S�֢#�P��$�F����I7�[؉���kRn��T ]K��B�0��)��Ϣ_��~�W�&#+[}#�x���W7����ܜ�㇡ [ ?ֶ9��%�ݷ��[ODT��Je�H������7á�s�%V����E��K=�j*�g�5	ߜ
��)�����S9��񥠷��1|��p�����En��(����l	�硟�F��o�O�N��~7}�&yA@�3^�����4�郞P��p��Y9�GzzP���+.~���}����nk�W_�N��?B��;���߂�j>G�W�Cy�̟�_���d-uX1��`��{\��c�Ⱥ?/��g!�|G:	�it����x�jq':��twÜ�L
k=oߞ. ����R��m=Z6�`w W8$��믥�(?��$��?���9Pp���H�����Ë?�$�+�nz�4o'����6hl[��itRˉV��0��̏�ƐY>���
-�N��+�d ++�Ld�s9}�tr����g��j?~�H�ƅ@z>g�v��u7V��(R��3ɲ��Yi$)L/��E�eu���B��'7�J���ݾ
0�]�k,$)O���8�v>�f�w��6a*2�f��t]���V"�	3�j������WǍU'Z�<�]���w�c��ٮ��5dP����P���f�z#�]���y������%�0�n�7b�_��+��U�6*:�/��i�f���O�A�������"\�Z�ZI6]�������f��~E
9/����(��+n�*w� �.Xh�DA�w0�{���������k�BQ����[���w�.޳{+���j��<Ǟ�W;t���)��]�#���	�X������W�It����`��YOC�(���#TI�?��;������3*���q��b$�`D�
R,�:D%*��P�m�Q z���Hs�л�J���;�����?�g09��}�^{�s��y����0��R��.���C�:F���ky,���������|ӫ�7l���,�����j#���8��������}J`!� ��n�$�j���״2)�d��-������6����B(��^\��ҵ&(��Tjj�M�;� �4 £ҕ�c���>�{��F;��(P�]�����VƦ�1�Abo�>�R7���cUzi�b������9�)DB�lQ_��H%�F��vU;�؅?��c�ޑid5|�ԑ��^ �U��DD��9G���UxJ=K�LG�`����x3W�L]/��$.]1��	õY��\��'��#F0�W�2[����p7��ύ~�*��K,U2}�����f��X�2���=Dz@&��<��~u�+X�/�X��í�?ݏi�K`��B�NrC?�@����"lM��o#����HD��#�������^���u}�k�\�����U,������qo
�ajS�𠻰���Ti$�"�f<�a�:��@e:v2|�3�;Us��~MSǪP6��4|�)/��A+sC�r��ז.X~ìO��y�s��������:X�Gw�ݸ�gJ��߲�v�A�!���]\$X�ښL���^\��������V�ӳW�nmc�]G�dcx�V��qǐt����"��r�)�{����~���*��5��D���]E�WݣY�n!���Q�W-�M������W��pa0�SS���;`zƟ��2�o��ߑV��W�z�a���T�4��Y�T�<�#e#'��*w���"�տ��0,�������M�>�)�ǋi�88�ﮘX����M��M�R �"m!=B�B鯖HJJ��vbo�������3�F\9]�1�뵫�M��(b���/� �7����w
< d�.;�=n�C=O"�-0�O�>}��ԩ�=d�-˔V(T�=(�"\s��Ks���Ay155ݷ�$���gμr[��ҥIKό ���c�u)))V|��b��S@���~�$�Y�Q	A�zf�ŵ�o���*Ў.�D/�?�8$*���,)E|�
�J�N�j�8��ޠ�"�%j�o����ɀ2�crL�����P��W��\	�>	�s��b(���F��u��n�惂����o�cg'���@������R�377Ov��ɪH���}}��N�XD��?MN�r���-�z�������i��Sc�^(	.�[��@��I^ЀUJ��h����O�� i�~�wr>h1	�%+���+����y%���ϑxԝ�����[�`:�DB9��+ 
�Z�Y
���gd|Ϝ��V�<�нQ�Bi��ڃ��7���y+��.M����*����J��@7�>c�&�[{Ztq��?u��������Ҳ��vHW6����廒LW7w%e����R��n�tO�����`��C`�9.Ns?��H�l�"i��>�N����)C+�O����'��p�e��_��*GRx3�LPV�}��Ý0�1����
�s��� �����dg��ݩ���^�Cȯ���6l�I�;c�+��lI���*a=�N����J&&���]���~�p��!�z|k۝�c̕CX�L�^�U�g���ݲ
���xiD��Y1Z�330S]X�2��Q��C 9����lI��$#a%k *�c�)G��Pk���X%����=��=�$���T,@�.ɩ<A�c
���Yg�N'�|�u�i�r�#Rʀz>�17��y��n���!�qgT�ȄZ2�t7#q��{���qRx���-�/*?ӥʣ�	���9X�6qRH��tP�;�0�<h7n/����-�
�G���	'�	9�p�P��Jj�W>�xz=W.�tED,H��Y�q�b��}����b�P�i�A4��hP��)T �p�����b5.~[d��'*ߙ�� �^�-uv1\��A8��W�5o�ׂ���m��w�K>��z�ξ��*q� �mu+�����?�-N+�����t"5��=�/��իI��#\\]e��O-#s[�G���[�#rW�}T����{fN9�<���A�Ǧ�A��CQ3�֯�9Ԕ��k}6?feo/H���p�W�_�Fqt�fD��2�mԥ-MP 22k��A��6���"+�U��E��Q~������-��+SYiu�4���p�`:.�h(G�P:�	�LA�,��K��}�Ľ�����~w#���"MtoP.�ך�A���e�������swR�r�&VcS�ͅ��D��o�J��UP+a�,�X��2(���oܯ
�an��;=�h�(��t�)�g����H�d�SיA.�G��B���Y}dsp�3���%y�Pڃ�1ꀥ�� �p��!ٷ�K�� ��``�Q�bf=�2Ҕx���=�s1���T�.�@Մ2�%�,�x�QX�B�~	?z�J\�k_<Ճ[��(��[L�[��F�aѭsHˈ�sP\5��ǜz�p21ȡ��9A�b��t0w�ӳ�C�Df�E_g��c��k�!��E�E�KVR(��#sT��qJ�&���؈�׷��ݭV`e΀�;���N��"�yx���_��\q���gE�B����RЮS���@Xk!����P��;��+?ruq	�Qq��(�Mp��
3�+6j�#�(L��y��́��Nl*�^�?ѿ QΗ�M�v'�Հ��;/b˄?]��Ugg�]�N-<��z`~�԰P#�0��6�:_�)�Q�~�������PYJ��V��ҢV⤶H` y�[L�4�Gb|V�튟�Ӆn������Q�n禉����حx�9�L�s[�\dPQ�" 4JEK&rm!o��%<������-_?|��<տʠ�U��'�k��D�i��`�@qa��͟�i�œ�|M2V�P��/_�y�HF��������V&J�֚͛��MO|t;�#�D����#Em��+��]8��>pu�z����YD�Z�B���AF�q?ݒ�ϫ5�4��$��`rې�6ʲ�������]��E��p��l>��9uK!�Y���nNؾ�DDF.��\�(��t���1��Y��>J7�j*�`O�qxOq���2�S��sH�t#���Ur3X�;H� M�����
�!:o!��zᎺ(��	��'��׽��e�Ց���+A�?�,�YL!>��E��Q���[�f����XƁl=乸0?�!��["L����9��
nU ډ��a�/]�7Q����<��#B�ŝT��ݭ@�aK�/1v��sBQT*�B����q��lE?�F677w��_�o!�$m�bR��l�����q�Peb��~���G�Sp����l%.u]�L��xV/���2�{va���Bw&�9���-�\�H3�W�\������j��r��rBI���}�s�a��`�Iz��b �'���u��x�>Q���Ah=
����~�/OED��mp%��B�b����� �ٜ l�Y�d��+��zq�ዎ<��i�F���#�J�/eD�<��u0���2�'�!�@�^������c�ߑ������@��� D����Gc�q2�ᇴ�R��f���>4X����H�
�L����84�xҭz5��/$Ǣ7{�Om?��7r���;���8��w�D�{<��a�����	��W!���G+3��H���wK��RV�1I�ktD�97b�b@s�]_�G���Q����Ã̺��j�F�P��BZE�7*W=�B�Ǭ)N�?@���}��?�)�MΝ�Y�J���8R#^@L~V�v��-��B@�I`�" z]X���m䠯���ᑴ-v~�i'qZ�K�a̡6~'�
��)u�3থ�H0a���������ƻ����N��ܿY�=����`SŲ`�6�`Sf�$i�@�L��{;c�̙ˎl���{�9+����?S4��]jb�y�:�ٯLԞ/���F�+�������b̽��Z�\��v��}��ǐUiK�A0l�/�����b�޺�#� <��HI�D�'��� ��@#��oذ!��O|BD�.��X��!��ax���ҫe�k��NT�ĳ�-�k����TD�2~��b�45�C'84��H�j�koޟ�M�ɾ���Q3��R��k��P�
�;w��"y��K� �y3�f8.}m?Z?���R:8t�)�b����ԩ���;帀WpS$4p@����Q$�zH�D�HPg���lGՔ���L�Up�9��߼��)o�53[Yh�9p����#*�þ��x�*n��x�������[A����Zg2��F�[��Z�WX�Ȁ�;N�LTS����S������n�'.fgAʩ�/��B����Fr���ғY�c�O��\�~����@��V��@�5Z�P_lf_f������"��>�s4�����,��b��\/��讞��7��/3RP8xA��'��͗�o���.E�ϻU���H�ə��[�j�6��*Q�įAߟm�u�*]>H|�L+��j[��3\z��z_�u)
���	|�o�mb�s��XM�D�W�E �o�+kL�EjQ�� �lg��DB�8�ĥɍ���W��[�8������w�|�<H����-A��/ޟ����f��}�^�j�S)�Y(Ҟ,����I��2����:���:�#���<���4l{
�Z6g�ե��F��4���9Ků��S�Ʋ�7�y�*{/xYz3%���d�v�\ڶ'�.�%��L���>�W�?�o���"���q��('�R��R����:i�Ny�ˑ�X�JH�\y�~	�ҔC����,�o~O�͛�e��d*\�#E;w�:��C���l�z�0�E��Yr��G?���s/�����ٗ��J&��Vimi�Nw*ؚ'`�I�q�z��fNyC�W�|��k�Xzۀ.0ǚ��D:t�P[�W�Vi�E���̝W��)B���r��tK΁8��
��Q#��>��N$��2;?����g�>�wV�Hv~$y�B��]sL�5+W��bs
��e�,����d~���y��n�}��9`G�O�����Qv�dXeE8C����9Yخ#C9���+�B{k���ve�4����H���:W�ƖmR��v"D��|� ��N~T�|VW���>����k<���" ڟual��`���K���Io~���_AE�Jy���&v(N�6��}� �nla��g!�9��<΢�jK���65���W��B�9��.7L�`N���xБ����f�z�4I�V=$͵�d�nٲe0�� V��8Ln��.�Q�x!����@v� -'�j�^^I��HM�Ӭυ�A�X��V�@�差_�fy�}��	�����4���B<
���Y�6��V�©��퐋���"f����Iĳ�ɝRi�ă�����r+�:�BCj�z� ������ۙ��:]�.�v��k�e߹
�G��=x�Ţ����������hH�^�r���NYM�)P��jjj�n0���06ȁ5�_pdO	V;~������k�l0�&C�T+�wD���Ź�s% ��3�M��Y��ѕX��q��q<k,M����S#����W<�H��
���899�:���V���=U��-F4�a�Y{�SJ�ɰ��d�(��т��10a�H�G C�����t�����y#��"Iu��vJ��יu�%~�R�>�������1�G����-�⣋��>��-��H���oϓdג�@=I�	_�t���c����dW�'�P�-f0��эFFF�o_Y[�	�{��	��W����o�&�Fn�:J~k���H3���� &&����R������z|��OTTT�����x��iJ�o�ߪ<������q�9'��w�5L��=��^�4ʣ
H�-B����� ��(x�l�Pd�*-Z��'�8 �r��k�q{�����ǂ�u�=m������lF-�ug�?���c�P���{�!�s�ls������΅�~F�%rKxIz��2���6Ah��ܽ{7�h\@I{+j��y���(L^Ԉ�����=�9�!Y�"��)(k�OTtڮ�^e�)�j(�<��j��g�� �(�>�Xg��������ϯ���y�Ef'�a��=UB#6�nejC�z7�xw5�U�Ԓ[Ԓ�\³_!xC�F �U�sWQK�c�''8�w��� z,��ݻz�p�GORQ"�΀��~�MO�
�ȸͪb���7�GH!I������i��H��˅_y�-oy��ŋ��'�}��(�Y}�����+p� �%��&��/���"҈R��ACVFƧ�0�k8_.���ԝx�@س��@��SVV�-.����p�z����%���9F�ra~�H���)�J�/�U�ǏȖ$N�����SE��mXG��:�sZ����>on���Qp����T� �`�o�cb4)�|�f5Qw8T,�3�N������7W53;{��VVtK��@����Ç�]'[���l:�$�E~��`��~�t�20~2��� dIz�Y��*�w@�Uz%rXU,�皮^�:���aD��8�ڔL�U�q�ι��**+@�?�D��-Y�e$����ŝ��X�ɭ�C@�� B����;a0����c��¢/T�Z���{��{(Q�8<�����>����S�u�n-�[��;|xD��L��m��960h������f}��Z]6�s�H�ZZj)��~!o~6k?J�_`�oB袓y�^?:kTI�������&$$�F
qe�Ls�^]�(���R
�˼��p��;lJ�F�ts�%���탨v�ƞL#�Pu@���Sq)@�u�QXױ���+{	ն
�&�;�gp����JX�d��jn�8��W�\er���C��gv �KG\ߣ9R����fef�g@~f֍��ui��|�(�q�R?uE�p������P�+I� G���e��?�u�+^�vS�Z3�f��EGvk��J3ss�u�W6s�?�I��a�]A��9�D<���{�QX�n���_�par��<a�S���؈�
J�Y6"ۺ]Լ�Z�b(HzU��{4WX�N�j	w����b���$s���1	���̤�Rc������>��kI���¿��N�i-7����jr"�]SOoo���c�Ќ��4��A.D>�2��+k�2Q�����W��W\]��^l�pΔ�j���m�B�*�H�r[|s>db":5�y5p�q�)l�H6F�w�&������?K,������vbJ[Z�Y���k/�/A7�r��7�ڜ�����H�����ȝ��34��s��d��Yii���N���V��<��迁��v�'��?t�8�#!�3�M�J\􃃅��5��wC�[[a:Lօ4R���]�v�v���fسP��k��L��A�Uk�Xx�I��D��ߑQcH�
<e�4��i�N!�z���~<�c�#lX�b�L'�����{���x���J���ѳ��+�S-�d+�xeK��,2�9��N��6o�s�
����_+�p��������4R�[���ڷg��95{f��\r��N
�<\��?z(ܶ={���z/����q��azO�n�h]V���6�P777�?5���GVn�̔�~x�ɨ��x�[#���B��Ke`��wp�����C)�%��Z#����N %�3��~m�ǉ^��)��eo���4�^zr��=e|��5��|�̠�FJ,�]�"�C5���}�5�5K0b��)6^� ��<��;(��7��ٙQ]����jei����m�sPw)K��É�7����QS�l�'q"���xfI5M���������o�)�E�`XeX�0H)�~�шς��;e�e(�f�f��=j�Z��o �wv)*j+��,�yL�v2��u�=j��4
C��7�*CҎ���U����w=OJ�;�3�GCB
g���}�˪i���ϵ��4��ݓ�	��U�}�|M�B�K�"��I�A���,1n&��KSs�_� �D��so�M@�CUcd��ۣ��Z�Kh���,Z�Y�`ӹ/�q
5�D^���IYf�W�VU�ă���r�w%%%bԒK��3����a@�h�Z7/4�?dn���4���/�^�-Z�8�i+��~aFU��/Q������s�1�M �����pH5��)	'%%%14l�. �/tB��~ # �W"�P.(�(-�ZWo�%Z|��a�cPѢ�#ۭ0�������ΟE���[%D�{�RtvJ���-B{��}�����s&N�lR��f���Vj#�	@�
�fJt�_��^b�������f����YR���5t�Dx��RT(_Sab0͆"�G)Z),�!܌c�?=[o�[x^�u���9G����.�����ɇ�_�\�3����2��Ȩ��#��v*��h�0켬�c�5����i>��2r���������O~<ofW���}�{���;w�.y�!/ό�p�����>Q8Fr���x�|$\�|S��qJα� �� ;�U뭕��Y���Jy�_��Z&��[?ۀ��!man�o�m��`���tFx�c���l1L��_'�O|�	��iד�&�}pҗ@�*��@���KA�xG��ߔ4r(yG�^�U�tyB�5.7Vkfe�>�oE-��������"<}�c��&�Xli�낧7�[���2)�@���Osdg�}e�ы���4`)EZ��o����8?Yt�̙3&�T��1�vM�g�X��5[�ju�zw�(�xFE�%��Ve@9b����z�/�0��5�4WOF>����ҁE�%�VV51;O�
��B�޺�ufVP�3^�L�7���_��whRL��V�jx>E�EX�#Ti)�*��;��N�LKm�T�p>$�%��C<++ַ�>�SL��P�b>����گ\��!�.�[�*�k�+���Cp���dKMɰV̸�hW����
o*��ܙS��!����ВZ�X��7?nK�G�Lbxl����F�����ʬ|gf�(A&w��������'��h��=�[z��<��)|��ķ39o0�:�wԍ��/�V�ރ��-ya�{��9��+k�}����F"!#��̬<�=K,l��3�+H'���Ƃ�2��ԅOh��u	#�{y+��I�s^d����p��
�z�>�!��������)�S�sG��>�#:_ݙ��=�n�@��S�O��.��w��.1�H}B���K���dwi�t�G=���R�=�2��ߣ�Y�:�%�I�rG��ϩ@�����n���
�?_��i����x�-^�沦��H{�����H��@����C!g�ܣU*���-���#FFE{�]��7����{@��.)t;`���+LB������-�WW
_�T$w@����/![�l)�&�|h�-�5����X���@ԋ���ڿd�׽�LI�I��$���>bae����a� ��w��2<|^c���/�"�oOe��6�y �-|�[�tch��S9s�?}biW�O-nPڭ��K�ܰ<T���EmE��A
p㊞���������=fS��\�5��͛�WVVN��z�(�+iDo;� �H:�$��^ā{������`V� ��`9�I6� a��:yN��K�jZ4��zlٲ�R��ij�cTԶxqDr�����7�.{���U���s�c�˨��sl 7.rw�S�x�:��8�O)<;n�<W�U����7z���(��Y*m�ӑ�f�F��i�&������\L��n��)�*�,�E�^�����&'�F`��_�::~�ĳ�,s�--AR�$��t6��� �X&��U��&���A�pHc��V<n�:tg�Lf�CF텀C*;�8�G��"��0��~M|�P	��v/�2{�9���G�S����)��}�;����NL�����΍���k���� ��9��ݷs�ab�y�
YVC����#���ꞟ�J�g�ey�
��y+t�g��h|/
���&����v�?�k999� ��X��V-g�͞��t�$�p�.BX=g���4R[-|E"�o�7�?���/�)7p����( ��4)g������� |@<��P���aNu�K���C!\�i�8���c��Ω_�N�XGj����߿';��J<R�eeY����y��hİ&��o�tD�E�@~�2��`Q���a+��<��1NNIY4��r#A���L��@9���Ņ{�Es}�J���9pOMm�x�$��$f)� o��U��dT����"������.Ϩ��}�D+�7�s��,�㩌����F m�SU�~��{�.��|��,��dl ��0�6J�1�B����O"��h�.�p
�,'!!a7���1�E���U��a1��㩙���D(9�ImCVp{�b�9��`��* ��U��!����۠��x)�-s8 �{<k�+��B��̢�9��ҫܞ踸��L|�g�tȯK�Q'���G���A�Y^'�����Mg������^���s���K4v�uh�>(��q�;?�{��P��.k B��L��*���~�u7�<C�}2ӹT��,Iz��ƨ��
�#�C
)���e���m�0O)�����5j�v9�LAV���9/=�mR��

*��_Ak�#�(�HIe,��*�(}�4�zʠ�!�a���%���d	��(>a������R�HX�SS���PRU�%̺"h�D�f���'�o�6�w�QƘ��0!�N�(O� �< �g虝:U�`�ߌ#{\���N�%�,�"��r/�@�R�h�`�|�{2�X��c,XS�t�s�-.DO�;�'s|I���R� tܣ�̂
 �~��N,�4� ���n<6Ч��
XCh��JRҊ����U#�rR����JBB�	�R����d��J/���������>9���O��**��Kn��g����h�~d���3����)!�	� ��f��T<�鐂"�mR`Z���o��EUYY��nI:L�����0Yqa�$����d.��j%q��Ϟ��T�fNX?E �@��9�Ü��[���d�W�iDR4$eE�.q�_0*�@α� �#S����A(,�Y`b,7���������W��=��	cc��(��(^n�w�N�,�d��R�Jͱro(hΙ��%r�S@3��\�R7��r<��!�I�Y̸�� ޓ&�ǣ����
9g'��ե[�IUx�;�h��tl�+z��|?�9T9���o������G2��QM�)�𰧳=J�	�A:}U�a�;�M��1|�K���Ӛk����! ��ng
ڇ���V�η���*t����}�R'xG�\ ,��Ϧc�H�^ ]f<�\+�`c�ԡ揢ʵ���]|0�+��k�����L���T�����z�q@�9f}�Ai����.s��(P�t���GЂ���
�)B�<Z.���L#���
�� ��Gm�)}@����g���C�B�� /��7v�oN&��#`�±3���x�5� dԤ���m��j���/R&��_<~p-E91��ehe}�F,��zR`O}Kۯ{��|�f�.�fzԞ4�o(��ʲ�����Rf��m�B��X�g�ղ���"�n5��|��Gd>�*����x�����Y��wk0�.Ő<.g��G���9�5DL.h|i�E'w%J���8�0�P��̶*��;F�����`�T��e�Nխ9���!uR����p{v�qʃ����F?(.:�b:�9�����Ox\�Sm�N��5��DR��^�{+E�<�)�ngx�H�����q��Cւ"b2�`�~m@v����` 'KK��ڧ�%�g'5r���Wlj+//|�����]�+a\i�/q���[QU���� ����.��8��y-���W''��~�^��w�<S�y�PGƕ[�/UE���O٫������z-���k���t�9��6��A|�I��-}���ؼ�� �x'+�X/������Wy���3���ٿ�	�KN���L��5���ݧ�cۈ����sf�%���#�W�f����*����jY��ޟ��6ĳ�ҥ�L��wk�B[Xs(t�u}ljI0�D{v@1�},&�.ށ��ؘ����b)&�A/XEYy�t��E��J�㧆f4�,K&�X3R)p�0ql�V6��nQxx6�l�{Q�"�7b���b	�`P���:�i�E��5�,|���Q��S��`��N&�g�aW�Л�(úXR8���s˸�e�*�z�X�p:ef������97�b[��fF�>����nQ�#�F�0z����G�B��ג���{�����@�تn��?>�τ�3 ���t
O��ܕh|�:[���	�a�ү�A#�����b>�� ���h��o�H�6Д5��i�D�C����篬S��>���%�
�s�����@b���������a�ٖ'P� ��$i$	�'k��⼖O�|a��/4�M��6��)��s/.�Xb�Lb�^I��r���A( �����hZ��w���;+7����Eu����V�4)y,Ϸ���?ȉ
6n���EN�Y�#$h�#�S�j�hB|��l�@s�ۻ��%ؽ-y�:���̩���(iikq'h@-Jt��тd�婫�ьAI%ef�LdL�����s�K��g����!o��3� �H��Z�>NG��K�r�}����u$�� ���K�"���x�'�zq�����das��uv�����, lL�ʫ��6I���9���ʝ�M��q����K?@�o����-�G��ts[L��I�ʥ�tFȧ�^1�"�5��Dfj4�.袸�dp_N}��I�ۣ�������sOI@6@15?�[R����'3��q�� �L~���*XU|�)�y�ש+ĥ�.s_��:�h��S�L4UՅ�=�ڵ{w�9�}���	ME��j A��c�ς��r4oSG-�ǧll�j+��r���(El`м	ŰWDN��_�~6
e�棸�B�Α*�S� ��`q���T$O�#	���d�&�J��kn�Gǽ���Ʀ�����z��\�hS=
���t3��;: W� ,�=�#خ��:H�������dţ/��r�{M��x+N@�XVS�{\D�	V��=�����W �U"/��i����P��0��5�$@tk�~���]�S��L|�W����C��~H����$�$���tzP�b�Y_��8��s0��x)|2T��/"�?���Z)[�"T/;�7T�[R��� ���ڊ�����I�0�{B"�%
� ���/�$-
+P�i��I�U!�V��[�v_�n�����E�4b���0^>�F���Y4M�K/kmՈ&}�x�F��fj�l �4��0�PT�]�3�e�O0�n��Z��^�k������#b�_��,��Sk��k���񙲳ˮ=w��HmR��h?�ܿ��j��9��,��X�&�kM��5�Uđ?466挴��]�ϔ�4ǐ�t��ݩsK$��W%PC-A����?�t�ډ(0�M �t�Xt@��ࢲ�e��w�Lr��ӫ
w�� 5�}�x���%�y�,)Z��q_=`jx�M<|����h#�2	�Gd� h�ªfu���KyV$�k"uS�mό���~���!���ٸ)�t�$�����]�R{�\(�9�g7XӘT���0E��%��w#��"u~�]�NԘ��/�!5y�+=��Y�B��=��>����p�wV.M<��q�Ƈ๹6��?��j�^G�k/����<�!����g|]X�}(����X�fX�qZn;����h�_��	JTp:������S��
�����a-ԇ�[�$�ǳ��ڂ�@ޣY�=�G^pT���,���32�onn�NC�pä��1����[�(�@\փ�ȼ�A~r��	�`l��!�M�b�L�C�̢�_%|�A�;��c!��oLTO܃Q��%��s؈�Vv����PKHH�c��V�);ҥ����f��o�m���$�m�}�&��#i�{ >P��c֓��	�A.\7���5�My���ߢ�E�fɣ݈Vbx�S Z3��T��܃�0V6�5̄��n�{���D��`�|g���*���Vui��e]^��`����.v�.�� 8����~ma��u�gsxC�x�����?�[���D�0�q��K#m7���o��MU% ��%��c;� :�*�7㓹�!�M��S�KhB��r-��G���m�Q���Z(	|A���B�_�x�Ҟ=g�u=�w�~�q[p����e�A�I�d��(���]�f�3�#዗��y5b���|+6���	�`:��	����7�.ҎgD*� q�UZ�i���@6^��/y�Y#�Wrh���p
��.$�D�Yӽ�e����&����jʿ��>�@��T:]p�p_w-�k/��8�T ����7v��*op�ie���d#C�*j+J��\���̬qbg��{C��a�z��Y+ۆ�����W���_:����&I�.P��٠j�I#mi �5������u�W0(�즁������ S]F�u���aށ�P�7���M�2�fp��|v+i4T���_n7��,�%@1��4��~tRKe�U�8BX[��]�z�����`��W��:Tql�Yƽ�(vg4����/�=�,Z-��}�<�7?HDμ�ęn�]	{%����NT.�:>��n���
 �5W�Q�
X��1x��"m�tR�ޟNݗ^J��F��:%V�֬L���]d��Ɨph�-e�"�����BS�"�Є��e�ӌge9rd�R�ްY����c�@�񰥴@��(��x�/�9�S��uK�@� �V�����0����r�䨷�,��b��9��V�KGj�&M�; k��ޡ�܄5��4�L`y.�g������5�#�
��i�7���"���*M��̗�5�6g��UV����`��`��4���N:@�A��꥗
����H,��(�B�ep�.x��>����Q���< ���'�׊N��YM�B|. �k[*$-�^���!�ה_�T[w]���s	��J�ε�7�.lx� *`�	�o�͖y�2�r�(
n��߯�o���W fd�//���Z�>~ l�>���䡴o9#�{�JHƕK�b	`�b?=o�>����������ט�6�v�_�:$�.;��o<(�7�)�R[2GP�!�ve׮]��`v��Y��x:��?�fo�i��h�4�>;o�W����9�H� y�2)�ݣ�] ګ��]'qZ�A����g��7���nm�@��H{�.���ێ;]<$��
^��y
Ի���0=�ӧN�`w"6?����~���7a��Z�!�k��Am�knL`u6@��şf9�J�,�7S�P��L+3�N��  J��E��]�i�y��#����:�ېbd�eT�6�$L���W@�d~]���1�u�M$,փ���WL��R�>��� ��v
z3��ZT����� QkVT�6T$O���n��˂����N�(#"wVL�{S1(�y���P%�G�ȝz���=0m����rg&��_�TO�ih�ȟQ��@��:W�e �$O?l!��A�*��'��c��+&��n�=sb�.ŵ���:ŝ;�ԁ�
B/�M���-�͸���DV�\�>O�,s�Z��,,ۭ�.��V�������ǆ`5�~�^����?�
Em�w�}����Fl����V�twd00�#�-��	-o�2(��IfN=f���H���Wk���C��\U~æY� r�:�j2�Ж���QlBb�Í$����L�0��7��Of������f�����f]�%�z���Zɕ��F>z�����]��P�1ŬO�a�N^��S�4)��u���K#_Y4K�)u���8$�{�~	�Çm {�a�EDD�yx5/dc�j��V�1�?� �J�o���oM�;KD���2�t�? ��H��y��/`sh������b���U�c+hk��)t{&�NT��ei��5��%`�D�oq�Q>��	}b �L�%A�BEr+�s��sQ`B��oa��p/R���KirH!&�����CP���F�d}PC��,��[+�7��J����&���.AA���8�K,��]��,����A����cɂp���x�V�G��C�%��a���c3�-&�Q;�w|�<�s±�pl|�6�O��$b��>��d�U�����^�/�zN���������+��e��Xn�\�M��S񬷠�M���p/�h�]���|����Ӛ��91�?��ı��7��O&O����M��
�1��aU���y���s�c������nb��b�t��w��HUo�歼w;��I]���/;��eܾ]oZ���s�w�p�>�C���O�^�����o޴�CeO���n�d_�H�8�b�:?���V��-X��S�7@�%�>�M۞�ֱ�e.�m"�ᮈ/'3}F:M.�U`���R�gs�@�ۇV\�o}}�O��]-�4Oܳ;F��[�Ө�-Ļ7�iI�Z-!b�T�N���L��Ů����M5;Sz�t�C��e�">kF������?���P�����^0������s˳���1��ؽ��� A|��g���ބ�>(�z�d�V����t?�i�E0,�^�:��SQ�
�^A���Ù^���6��-=-�cm[�� �W=R��G.5QR%��ߛ <=2����k��s��m�j�M�}ὒشѿ¹vxx8�/���^ۺ�0xsySv9e1�5c�֓]���0oAb.S=<lH��ɢ�-��!������?@E���;/_�\{y�u�(��9��/Z&��T�t�=s�E�i3�q^�zzz���C �nO�.J0D~z;2��C�s4���[9�Gj�?�QV�k��"�Ж=jh�����w��WX��k�k�XBػ��6�K�XX�#��r鮲@Fҝ;w��lR?Dus�������NP���%w����VP@����JS���/D�ʱZM��I�#�t��8fM�%���j��0��1�+SQ�:�q麼���]����Ճm�ɔ�y�yU�"�L����'gm{}`=����:��< %!�s���2���9���51;�E�q�g�啾}��n�[���b���p�l�svt�6�J"��}*7���B�>D��Snl!��k�W����;�ֱ��7)��cK�G�����7�ƒ�H��*�!�~?@T7�ڦ\�򩄬��q��wY��6��yDj��M�{�tc؊���=$��� ����py�l�0>�%�ܜ�ajbR�Q�O��Du�������`���M*�"Xe-X�Ӽ���O}�����!��\m�xE��[�wL���gߒGFF�
̉G����$�J�MNN>�:[�Ј�߲^���c��?�-'d+���ӯV%7.���Lp_?y��R��q��Zi��g�
A��K�u��l>g��;���&�
!�\.oR/0Nj�1{��>	1����"!z8�&�.���mdT���D���L+�L�y.�;`P�]�m-荣�?~��v@*K�#L�v�)�w���I��7Щ���+B�g���Ͽ����YQ~�F��9�!��TW9��{����Ǉ���zk���\.�eO;�yYA��>#n�)3��v��V��{IO�5��JNuɱ��ȴ�e�+.+w�[�Vg������.f2��\���i����)�A������@�q|��u5������q��J�٥�	�s'tM��^��]�X#���7?���������I?Z�E��d���D�,��9[�O��A�%���F�Qä��ߩ���!��#��I��?ݹG~=`X��F�Q��4�����==�6!�k]��x7S`��u�VE+N^�VYuu��!��z�0-z�O��h�l��$�A���n�銻;�U�V���^��l0��u��]GZ��j�x��񔁡��C����'�7�o�8 @\ݓ> d�8��9ƉUF:��#�������7�5�A��U�&��[�Bg+�d��΃=�6$��@v7i{MQ�-8@�[G58b�_o��ؠu2vi��6�2W�X�Z�V���ӷg���L�!�˟n>N��j��O��>���h��J1G-��?u��ڮv�̔���q���;RK�d%�ٱ�x��lo����Z'5�F�`���w�h"�����^�¿�����3������mf}���3�q`�r1�����.('��D���FF!dϗ8��󙌜��u)V�B�~ġ�T�Z����q�1_pyjM#b���,���>D�9{��m]Y9�G��>fv����T��} s�i��{��AX-�hi-���������T0�%]�v���=�޵���&���WC���D8L���Ǐ���m!%�_se�����XTi��I��o���%EW�<�u�~�/�s�C���˿����U�X�����t�[� �nlkk��$*𤗖��â�;"K2u�m�s������V�� \�w0�&���������E�:Ւ�W�`
)jkL�ȣ��s�啊ʝ��?\����<DiUp�MÏ'j���]��'m�>}SM=���WR}�z~9}��ɍw+���i�E����c���W8s0�({�^� ��2M��A��
=z2�F�+�ܳo���Hɖ'���+y��XPD����@YY9��Nk��V�y]�@�1�+,�&ɔ/�N�?4I$4�5r��tχ���#C��d@�c��I�o�+��tA6�E�͇�� ֝* �v��z��w"�j��oj@�� �ͺ��Z 3�8�Z?*)������6���K��$��8Ć�>�����꟰����M�j�~>��9�<����Kpp���=w���a�N� �'����v?j7
W{<ٖ{�ں���q���Xn]ط�NI='�d�G��DqP��C��B2����!C!���2g,��%d��92��Z��y�������[���k�u��Z{�+A@�xR%��?�]�`u�ǘ
�7X$�d����
���O'�=�z��!����L:�؟�� gBJ'��qiw���h���q��0��}*ϐ�\�T��>�����P�ē�Z��Wl��w=�Y���G����������mov��D7:^k�p�>��&����۷������ g'r'w���eX��R����N��:	QS�l:g��W)C����bi�xV�;�E+��i�*�B���9�0�
�x׏���6��r<��A7
)�����d}���.��j0��������U2��z���7"��^pb2N�b[�����W��)3�p���V�W&�`�_@��	��S�����1�+���[��~�#��~��=,}���ӀN��4�Z�w��Bl������'�g�&���x��^�v6���#<ˊ�h����'��d��,TW�5�f�a�w�a���_ �5�lZ1}|����U��>`�Mr��)���! ����O�G�<�I�b����9F�%?^^�����67HE�����@��|V�f���M�z�� ��s�A�u�]?�gqq~]��`����}�n�$?������1��Q���[�n�h�+S\�Ad����f�hN�,|���	8��I�A���,9yd9$��">��/NVrF��9��,m��������M��"[~TLH���~b��k�#��J2�
(=.� �#k0���gr������f�<���H���F�ل0^��u�ͦ�j�,77W�d�/�$S�@:D�&��{EĆ�%��z�/���D������-!YVa�A���m`�Ǝ��n䔿��孉��ˀ{�U�KiԈſ�C�U�^�WX;���##�k��e�HfK�wm�/+�<9�'��I�&LD����֮g��c���Iɐ��ЀY��]���#i)�+�Y��,k�k{p![~Y�MI�"�-�0՟����O쑑)��kׇ1͕/V���%�L�x�p��8��o�."�z�࿻ �k�S��jp+��f�5��L�ԗ'�C�>�j���j����)h70<�[�Ա|ZQs��AR�{�to�WS)i���"E2&&&U�OL3��/�v~�3�"d�Q{%�՜��Z4GRu����ł�h�Jp*�3�#fN��m����
�	WI>T�ܝ����G��M^�65������Щ/ �a�k�s[����_�}3�Z,���b���˳
����5B����0A����}��C�i��]h�p�g�㲣]VD�vr��T�/9M�Y�'�J��zD��4�vPݿ�N���=��g��t�(���yyx ����/vPz����+����Ρ��l�,m�$�9w���?��*�Gs�Uh��HAof�U����?#;w��\[�r�ק���ι�M�"ۇ�&ơ�(����R�f����:m�r��־\Y���Z����&����MӦ��O�j�C�i)��z���f�A��}����4jPT�)��.0Okt �m���ѯ�|p/��!�|���
ܜ�WV-o�V%�j�YZckCC�=��I�_���|�m����&�r�=�C��p�Pb�"��vs�̝O,��~����S'a	?�A@X�죎E���/�=�?��T`�F���ԝH�3�#���y�?��1:�LW���}�	+��P@m�}�;9��=6��tkO����d�S�:�%A�ϫ��U����g)�pj���$�W�:��N����:D{!�q�P�=�i\T���3��������P�/�+VsA(W�څ��-<>�A���&������uB��o+G�7���z��=�G�9�0UHϱvEA1��zb�����N��^׽K"%`���>pްc@���٢�z�X�b�DD�\|���}(�C��D�/�m��`�ƪ"��W�����)Ym�F�>�A�r���Wp+����P{#�=��ǎ�kk�����}�/faz��5���v��!ٷĒ	ҕ�HZM/�/=6H)}c�Ƙ�B�$��_�`=�I�2x���e|��@R�y�_pu��ǖ�
UI�ohhK�z7�˅�1��JnZڠ=���E��n���ԕ{�/?9��#�*�	��N����<��2�T��&Ӏf ��x_�����h\����e���\ �q���N�5�b�q9��>1~�j��q�?�P��ZHW�<��o(�8z�Џ����Փx�B𢯯�,*�Ii�鑌�!$��k��W�\Gۀup�y���h\�X�/߾}��Y�JFk�~II�������R�VY=�Co���#�?O�f���Һ������:L^g!��H�%2G��?���ur5�RGW_3Ңq�"�k.Qg`|�x��umD����'/���f1z׾�U��]7���_3��H�p^;�,������\���NQ��m���d4UX����3 �"�lxx|��p����!��p||�K�˦'�4���
��)�R�T<���)��S�l*e`j,G{ڏ�'*�E����*ǯ� 'M�o��d�����ͽ�
�x:e[��X����{��b�~��$���f�{6�S��j�C���?v�B��,&Л������l����>�}q�S�D�\
P��,q×�#U��Hb0�/�!p�'I k#/�ՓA[\tֲ���Đ��D�~��������`);��2f���"�ի��J��{qe�R��Q���u`���lU�z��d�9�7�cY�(D���}��ڹZ4�pq�?�m�WJj�o��S+T|�u���vy�X�A����~���@�Q�|e***Y�����%�R��c�	o��T�~�z��C��,���"5A_�.!��Si����x�n�fi��X/��8+�����X���qn��R�Gaވ/zKhr�x�C5��q�uZ,��뙵lr���/;�܊�E
��,�߆q^mU.
YYUN�X&V(,��G)��n����+�J�e�r~�/�`�IQPbQ����~� Y�R�IF��	ׅ�Xb~�}�C�jw�n�6�.A��S�����Bʔ���@�_���ů�2z7Y���8�-sQz�A�a7��*������"u:�Id���O
�v��j��E�Y��^��� 9�?u����#�-��ªA1ovf��a�F�Vx�g�n��S�x⦖����Пl,���i>ߴB�MV'.�!)w�6�d+�����IX�����ԑzSJ# ���M�5�SX�||'�5l��NT+��db}�~�eF���˿���"�y��2�.��m��ͯ�ƀ�+�j�K��¦n�M=����b�f�����5Pߔ�
U���
���NcǾIi��Tj���Wǻ�3���ч���������W7B�� �R�%g E�Kv-��'y4CVc ٢/��r"=fi��:010�{�u��9j�oo.��cSʂ4�n\v_�6<<\�:掶�}�a bPhjj*�,4���R���ܛ=�<�1]��=z�g@���S��I�
��{�8�{q�5א�5-� ��}�S\��o�o�/	?--Ř�M�%%�Q���H�����0�B��"��ώ�������;����&WYBmw��P"��v��Wp@���8~	N��g:��D�ʗ�q�OW�Kv�.�7�%�l�x<�Zw�5��qU������v��n=F	
r�Վi���9I�'-���?��3JP��<�w���J��}e��gŨS̳��C�"���^'k3|L�M:�������h	[~��Ǧm�ݵ�F�%���� ݄`��������9���~�Z�oFne��<&&&�����zE+����r(M���i}��Z�g��CƓ�Ȉ`�����\��}`�M'?����j~��)&D�t��ӆ�_��D�q'�R������>؉���~��)���ȿ��~��R�O+Rw粣���=���?���B��9�<CZY��3f�� ��^����R2�[P"pj��ŒL$�}�A[��l#����b�����O�.�g�n����|�V�B�p��"��5R��r˔��&]ՠ"�N�/��}�'�"R��'�'�-����G��Y4�BD� Yw���)�'o�xE�]�O��v���]>��B�/V0�M\�'�2���������v4�v��:��mI�B$m9��R#�`�D���������Ќs+�#��?��
�W���R�ΐ�#��$�4�u�Lƣ�{���
x��/0��w�O�	{����-֣\,��>��˥��+�/yȼ>�i�����'k	�=�D8$�� �<��?2b
/� m5�jO<93���ۥ8�(U�/C"���C �%g�OC<�~�]�9��6��僫���mbA�|��l\\��ec9r��������d�1.C�ڪT?�G�#q����j����EX6�T���w�E�z�H��gj� )�|a�64�_�Ʊc�[����{^��O�I�e�Au3���9��eђ6���]���i��C"��	��ov���������ĉ����0@�/���9��X��*	"�P@��.���،��mJ>~�h@��V� S�~��-�]�#����+d»EП���F�ʛ�*�`r^u���2�췰8EۥZ3>�\� ȥ���p0ƿ�$���/^�5XBer �A��>,M{�V��]s(Y��`{/O��l����p���D�}����ܘ?�p�mP�٭T�� ��X
d��Z���P�2����P>�9Y{�!��y�M"W��Ī��n=�Erk����[3����}8�֨YW1hFqI%W��:zd	�O/'��}wV�Xl�D�	v�ky��Ƥ-�''�h��[T!���N>��8��T��@,�`-Ӈ�d����*!Z4��8q��vI�a���"�r��i������+�h v??�������'n���k�����W�g1B��U�D]�
���5_�}4
�&�(j�	.��oF�% ���7Q�D*�`��\s�N؁� 4�o�S:�y�?$ݬyn�T��Ȫrѯ��oԀ-Z�P�Cv��,�Q#�Շ��A2����ߓ��/;���`(��92�Ǔ���:����_2���r!M�W�ȟ�'�Jv������oEz�����<�ڸ�xb���---���:�A���O��K�Y�r7I�Ȅ
��η�9 ��Y��(D���$x� �u��^�C6��BpcS�(o�������i�ErN���j���/�}�ÎXˬ����NQ�%}�y�7i@��w_lC�!������m�ԝ��L�C�?7Q�$�M��w? �1��U���i�Z�O�flb�!	�����W��(,�\x���rk둶b�rϿ
�w._V���%�9�ޤ JMƳ ��)`<�#�����4"���M�Ż��?M�D�qƹ㦓oI>YĔ������6T�g�A��rL��0QG�1����@�~ʕ�@��t�d�`r�g.�&՚%Rճp�c⣷�w[��N�8P
�1#N�Kb43�dDD�qdR�N�J��o"T/�ju+|�G_�h�3K�	�Meo���̇�t����ӿ�M�����2%W\�W�%�l�o!{`
���Vm*��F�E��,��a{v�頵Dc�}����vL���x�OU��8	Nk
����W�ʝ�fiƓ�����2��E)�`L�X:^2|�lD*��a�v��w�~�B������L�&	��@���^�Uu��X�x�6�'�U�e�jPN-�cנѾHy�0��P�K�yNw�>�ڄw��꜁��nZ���PrX���4��	Ђ'j3�~������a��m� H�S���a3A%B
u�\]+������+�ݻ�S%���yZc�#�7͵�X����j&�����?u@Y[1|˧�<��jV7��d5����yŵ�:�p����VY=���Ո�wV����-�,�;B�|������ghu�I�kW���}� h��u�RGA�D0v���!))Wk�J��ܠ��U�A�i�k�ڋO>��?�K���kI'�=�-.���v�C���j���x��l�9�!����G=X%S��k���Q�����G�*�2�WT�D��>��n�U�����4�?���T��h��8I����Z/v
�Et��؞[�O�B]���/..އ-'���ߥN�E��[H����Vۏ\����t��> ���u$ٴs�h�Cd�y��'�`�T=�I4�Z��p-G�ip+A0�G�^�oZJ�I4H���%���X��,��;��K$p���Y�>0�̭]q��-oo�A`�Φ�x,�,��:y�ONS�Hlц/ҽu��������e��=�Ɋ�a�8���5�����c��:��79:	-�-��%���b[�|�]b���v7I�`��{�/�q�'�R)���������&�E�Y���:e�kk^0䛘a����	N��g�{j��1���[���~|����xx��뉈k�b���r������0~��_�_&��"�'7�;���-h�o������:��:�n9�S�[���_��C���}���:n�^ K�� ~�ۆB �C���VTD��O�TӮ"�X�\=R&��.6�:��&�i�+�
)�2~Ư*E/}Z����Z�&��u�Ux�5@yţ���o�_&pG�&�Pxx��@���@]��`k����sk	��|�j�Z
���ǇXɼfD����������]0/���$ԲӺ�3s����kؠn���Ǽ~�3�N�e{�����m��a;�t\�9_֚Yb-��hp.�S�X��4'V���y< ���;�y\��f�� z^��@����+�|�~� lF�������I��PXX�8I~ r�$%��,^�Yn�V�0Dsb�\\5�V���^�P��'s��Mh��-��W�!	l���^�,����-�۫������϶���g�4h����g	�`+��Z�@����D��;�v��yS�|xs���lњ�:�` ���6��SYYY����Q�-���.Q$�3.��x�g�b9���s`��F�oI���N�<���	�"��l�����t�����"�,�9�V*U�<��)�#^�'��2 eN��(�'O4�9���w?��]7�o�i���;E�G
���wp�2 ��g`�3�p�|8��R=f�1p9����2y���ר酸��0�<��B��|׆@�Ҁ�oI��O^?8��ԁ�6���_��2���Z�y�UJ��}׋���'6��ss�As��. )z�'�a7��l����r���DTl���x�!_J@k��c{�p�g+����x����
^<��h&���M�!/�>�`��������������ϊq��8����KG){?���0��� B�����L9l�6�����ː���s��ţ������f�F��}���t��Ej��Z�!��.�8�	�Yꚛ��FBq������B�Y�}>d������MB$�עiI$	�V&mݚS�t��N	��-�g��)���>�U�0�3�\�FS;��܈�����G��F1��ƊP�b����Z�ڍ�w,J�n�����V���d.Xf�Yy���䤧̀y��N|��'exI��6� ���g�>�w���P#�5#��0
g��d^;�n��G\��������
b�wq%/H�I���h�%�?�n��yL�L��_H�m��p ��m��!�as��N�p��|����y!�y���eMMMo�ƌ6X�i�D��
߼pߟ4XHkO�#`+w�3���`ӆ3����u�T�y�U75����m��;&��%[�J`���2��,5�-#�G��`�o�^Iޜ�����8�eJ�����R��D���������q�J�MUeew`2y66~D5膀�+Я�̃g^���v��>ò�J��!N�\�ܢĩ�̭��&���HQ���ލ������$�#:�\�U=c@��lւC�<��������'͡?w�ۣ�|w�QW����¦c��h����Z'�C�Q�O2On���0l��$�LS��5���/��թ�U~Z���C2%+� .�h}GXASb��n��H�K�&V�^>~�GGǬxO��$��c>;���� �czH5H޼�6ޛD�K��">
���%���Bo�H25��/+��^A^�>y�k�y��mvv��@k7�=d�
�&�r�ib~��R�F �O�D��]�ғ� ��e�@s�P&��Ģ���~iJ8^�������mƛv�W�^��w�2�D��UI�OL��Y퇻�o���ln2��0��������� !�$����+ �8���[U�nW�MR�Q�VV��w�
��"T���p��BZhH`Y{=���y�aGN:x3������&ĐΜ����*N^�%�(��rf(�3�(fIh��7YR�o!�0M��,�u,�i=�/��E�l�����?).�d��@;���'�i��%�������Z�k��1�w�h�B���mҞ��\%��l�?��M qȌ vpQoR���|de�^ԋ�9sbU�Γ(��E9OӺٙZF~�U��ׁ���߿�F���/h�����4���
�gX�W���$1�uݭW�澞��qxƼD*�ҥ��:��u�2��:��;��W��7���]�(�LD�}�c�����+�%������͜��Vŵ�1L_�=�J�h�ecFj�~,��~t�ݹ��ˎ�����ʃg�Z�k>|zy��q!��{x�\�Ĭ����Ȇ�j�@�y�������vhǽ�U�V��г�eG)����>魪�;���`�ׁ��R.��L�`�X��,�#�[�>.����B�QR��V]]M���b	��{ʪ��0����HPw���n�jx���@^O2�;x���{�k7?��#��g��%������Q�>x�h]l|�F�8Ԕ�^����N�k�qgf�VHp�]�'�<)�̬>Қ;�K�ACC�C�扩Gj=6#8	LO��v"~8{sx%�Q���{PU���;��)�Ma?��'��N��FX	H���.C�4�	Ss���;�4}����+(Y���Z7+�A�����/0������ZY��;�4o!��gw-�v�]
z����9�tH�;"Ov�,a�ٲ���������6�~�lo\���'���o��j$�����<����\��)�� ��f����.>�>v�M��)81Ծ��C[U��OW�C�Y#Ng7T�ՙ��F��3�l[���>����#^�T=��74T�����`p�����p[��oʡ���WGX88L�ad�
>jYV�l6jǎG(��w�u��F��>��  �xȑ�P�>Ԕ�d�ϗ����E�|��'��¾$S;/SF?㯡V����z�����ޘY������?v�&��'�^����{%�����W���]Ğ���#��V(�/�j,/��N�^�nY�\�u����b��^�nm+�k=^F�n[��|g����of������r��r�/+��E���FB�Z������MC���ƴ��*"�{ӆ�����[%m�5��sy�S=7e��+N��|;��H,�~�������xl2�lp�5.�sv5��M�O�z#L���59�&��(�<�~�ݑ������q�_�#{j�X��(�l�*����̮�e����-��ؕ7ݙ�pV�_����kXM�GݻwO1�B��m����%)�\�lV|8_�w���_䕏I���s��[����T ���o����e뺊���HN0��B�,Qw��_��a������1s���7]�z�񊲕#�.��?��C�>��D�M�R�-vN���a,Wsݦ8Fx���-�݆j.-�R�"C��U9������~�]2�E��ǈ�LL�H�ѧ��}���i��2�4�#���(��WQQq�.|`���Q���q�ĬW�2i:�Mg��j��l[K���b1��1�����ѼJ7�u]Mߕ��\�Tt��-|�C~�.�����gg��M)���������
��[%l�O�B���a�P֔�CN�L��c��.x֡V{e4��^���FMԚ�-�C��3�g`5�\��sqɂ!�n.���`@ۗ���K�/��N��l�x:�bƏ1=K�$9l��/ W�r���Tw�wH.e���ϡ�T�m֠������Ne�=�xt����:|��ޣ����ɳ,;�:ɪ���M�����EF}�1��Â��)�D��v;��$�X�������LVuZ\ͨA��2䨨i�C�/+�p/Ӑi����V�Ǎ�ljMsw��F|���+��-��s�%'bh�`@r�A��T˒�f1]����Nw͝���ˇQ��'�h�Vv�8�:r�o�!����H�6���.����>I�8�������*]��8���w94�*�.E]<FFb��( � gr�Hc�s��f:��"������w8�$TKC�?��,��f��1�i���܂p� !�;�X���;V�ׁ1���sn�b�:~���q��L�f	s�����62��_N�,�KV�?��֡��B��<i�/}WHTRI�hg�=�W���~�~�~_�@��S0R`YJQ��D�gyO{�E9����h��p�������"�rQ=�dG���_�0at�_�}z�����Mn�.��@uR)RF@����J®��S��db7�\kў[g%|"��ua~~��N���b7c�I�tU�G����&�E�����Z���I| @"�2���u0�S_Y�E�]���ٴ�����a���(���|A�r5�6���r���F}�b1��w����E{ى0e�>
���}I�O�v�vj�m����m�1h	�����Բ��?��fі���p�g�`�nff��/�����¢;�a�6�ք�V��7ׂ�}>i�?���ĝ�M�p�؞�A��;L�'�e�v�)#H�>Z���7�iu�veb 0� ElS)
'_�M�X8B��﵅jU�z\��3�&�� e�(��PN����
�+��Я�S�f^�Z���?��mdʺ
̒�b��������O�T:��"{��jj���#w�ү3{y���V9�5����Pϰ.�V�� ǇZ�~�j�G���5�، 0[��;���u�k�����j���M�X9�P�	 j��x=<'���o&�`�<�����R�4�M)��CGD�(�͆�*��
�:�4>��c�GǏ����>��|ט�˻��0�G������>�rգ��a����#N�z�~��mD�H��֣H��D�At��Y�X��V-��`���C�փW�U�� �������y��p�>�6l+���7$��{�&@J^���ħ)��9i�P++��k��BZ	>��j�O�= ^}�i㥈3U�A���e yA��q6o�r	�gN�
�S(����i�:���)�����*�ÊȘ�h�^&�1�s�zdC�"���(i����2�q�c�����q5� �؜I|�����e�����e�")�8��V�ЯN_q�2.�h=��^墍��g�G��)��c�eb�ూϦ�߀�<�kj�T��S�%?7�8<r�q5g���Ϧ_�W��5��hr�"�c���$��W�yt' L1�=�>�����ؠ\D��������o�6E\�K���[4�� [��Us�����b���c�D��i�A�	e�S>EX< &0˘�ĘyP8~mpE�����ٯۛ%r?A��>�u����m��w큔ѻ�Ad�5A�F_0/��x�Ӿ6�
�L)�@����v��
"ux9�vƞ������K.�����.]_���jY���JLvJ��*��|c*-�D?�/&�n��q�E	�8|�:�u���4�pK7�.U�"sQ�PZ�P�7�"�Y��?�oW���]Yb8��+O�rl[+`B}Ssq*E|ضH��ӝ&q;;0�P���'Z�2$�'!aB>��2T�5��&�����U%�;M���߭W6~,��{�v��|�+[�\�Ӭ�,ZQ�r��d��˷�(4�[����~���@͆���Y�~��x�/0�����ö���B �q���JH�A(��3�X�G��[?�|��,e���CO���t��a�`U��o��D/�����
X:�ġuBZ���gr���ޅVK��É�]�!8� v����죪!������.j'�a��6�J�4���!���늚h�F�����V������|�k*)9����i�~d*��z\��tV���&
�gi/M�׋m%��u&�ieW�� 	�k\�M�}X��*+G�CC��fE��\J���i�tqll��>��l��X&��#�M����N����n�]`��&.�i��:�F6��=�aq�`(� ����<n�`�RB���Ԝ�#�M7ɷ���s�|ku�o��_��� * v��ady��ի�K�奁���P\o,C$��8w���M7�	�e4��h���T�,��{/?�x=De���x��={'��
���*_/�_D�������^�$;�5᚛�U?���q�k���|� �7S0_i�M��r|m�'��n��ی8|��v!�lv�6�'��+%(iu&&2����;����+��#|���:�72�1�惼��!��6~��C��-[bˏ+��_U�	 ��� �餴N�49�pLr)�U���G������>j�/����ߨ�`������~�q|���#G�(^�?
~t�� ���ھM`p��0a�L�_:��U�i��i���7�F�L���#���!����և�ԨMa'�݂5Ƹ+�r�U�/�ؘ<�� �f5�,Z{Yp��P�P�|��&�
�9�ǩ^<Ŕp����G�JSJ�&��9�2Lp�p�M��Ʃʪ*C�R/�+���h�H�6nʰ^��Ǯ9�W���{I�(��i���t�Ѷ�hz0���P��W�[���<;`�𙷂|]�,	�~����.�5g�2�5��P���h_���n1>�|��� `�W�����J�qW�	�#�3??�n6�)��
�Crc�b<l�CvK}�~��Q;�0�H�t,xʏ���ه�.�M)�(��g����n���$�֘��/S���X@(577��HU3�#����	��l߄�5 �9�O�[��|�R���' ��������f�ܺ7a�� �
 ���Sǔ������+�n���FpƏ�V}��KA��荫r�1u�y���m�*ii�	�R�����a!�3l��2	D0>n|R`������Ν��W�:�ດV�������&�Y~���2<�\ĳ�4�3���� �as����p����9��f<�0q�����VxI��v�Q���?A($�x�'��94M5E���S��Ņ��^r*���ы�:*����Egps����u�@���!Q�ᆻ���eg)P�,uC,��"J���)�w/�߾um�O���G���jcZݟ�^&l�����1Q���*J>�F��T(�r�ۯ���m������=t�	x	S��W�o�`�8_��Eķ��;[Y߂��^�MEӦ��� ʘ���O�1k+�X���=>�hB{Z^t7�����gWs����Ǌ/��#��3C��CY�I�#���Sy�V�M�6�_K%����'y��5�f��۰�)�a!2�2	'ky����[��t���8�]���X���H�n�M�+yY���R����>\QQ���L�+{A/���<A7��/�*��/�^�;qiiqa�hl�.�w|$�2�d�ˣq��p)�JD�!�<����L���5�����/,@>�n��*ڳ���qż���_B�[3>�ؐ�K�˴����tt�����u�#�o�b;�a�`q���M���O�-X6l�i�r�3�~n(#+UWUҊ#��u������X
8�""�Nоb^5Q|:���V�eZ]��M#G�y>�9 ���GE�o��a)m'�c��cX5����-�c!��Nq���Dy�I��t�ޅÃ\	�� 	�}G�g��dAn �s �8�ƺ���L+`L��]�j��PjM%��ĥn.�_I<��Ue�NZ�&&��IX��3�Y:2k�+���Ha��S�'X�h�� 8F]�gS\�p��q���P[h[P�����Y��[��,�8�O�.��]�Q	P�Е: B?�a�-�N)����5
FO���t1����ծ�4 l��? ��)(>�)�"/ʷ�"�m�~�=<*jɏ��/9uV� ����n�*�6?�-�oct��݋mv9��U0���2e�<Ho�X.������!Al���q�F׻D�+D�Z$zp�$�	`�U x�qc
�]��� �mA,(��aGj-���NFԏ]�kY���v�Z<ʬ�/�!L������I���X\y%vL.&ڟ���wnr�͈&���?<`8ܚ;W�Zp�)˾�3��4Fٱ���	��]�b �������w����[���H�<&�3�Vg��Q�oBM�����	�r�����Q=7��<熰#j�1�l.VA�+:��XC��.���,����㊡s해�ʺ��^{ѯ�����j�f�¸cd��s�!�p�����S;v��y>�*��<�������Ç�<_����绐});_�T�B�ی�W�3��ʞ{Z�*<��u?��W������ RC��+je��j�I4��U�|sd�}G-���{�yx�џ���m
2X�M�I��*|\��p�}�">�mJA_EN�%°��zsG����X�(|���	8��ESim�z6�5X�?~ �x��H�	�h��`�Ƣ��F*�~{�='�8+&��׻�I���L��Wӗ�	�Z��8����;�n���D�0����(�$F�m>��ӄT��V�����+�l�.c=�\W���݋*�g`j>�w(�װ���hϚ#�����cT��Df�S�/,D��
�X`�"�*x���tDR��� �V���=:�梇]�F�>���aw�v�2�#b0�-�5mޞt��D�vt���6�ߔG���* G�j̰nӭ���oZ�w�����q�M�����L�q�6 �K2�]����XW��\�A�V��hʕƽ�t_ y�uoc�ꝇK,�09<�*P�d�S�&U`z����i�LH������lp�8�������#I��Ċu�/��
a�BT��O;���8�¹�*{���|���rd ,���	9l�EH�|֞����-�9_��T�<s�XMMĆl8\��l�SoI�6rdP�n��*hᡀ ��v�Lh[K��\��	��1�0�|G���2�]埜 ����\Βd��L%k.:��߀�h��MBB{���C������v��6���Td��$��z�]6��9)�� R�-�J�~\auU.�b[�ǚ�i�Z�rL�g�P$�\��`�awk�qv�o�;���<�_�v��=����D�W}7O��l/�:w�[���y�e0s0�(�Ѥy���H�,�S�N���U�f�Ȯ0+�_�8qcچD	��=�i�A���hχs8��{wI�an����("X��qs;�pO2����4�h
��bBڣ��a?8]�)!�w����NV���R���6R ~�)�P�����L{-�����Dw`����@�d�fn��#+}=��¯����װ���涚��������[��o��4`��:l�E{�)�2u�L��\�@XF����ͨ����v���L%c�
������4�ه���3|��&y%?WU%׹I�L��òC?(�m`��Z�������*El �
4i�}k�u�oba�[�b�8R=O��`��U�!#�[/;�1�-!�Wq�K��!���a&��d:���g�@�R��<�j�i����b���Ķ8�a>�=OeG��]��\�������	�Fhh��f96�٧�P�ſ)��_3Y�r��4�WLU$$$�`VK奫RT�3��(���}�n�%'	9p�]��9�H��7
"+�����إ�ļ�f#ѻ�`��iE�R�G9yAEQ��񌦅�� ���-�)�� ������'�tu�:���YGi���a�ػKLl���4���[X����-���c�G����v�%�!�<;\�rj�
"�3�E{(�b͹Z�]��a2�%>Tb��w��	���7F�-ڹ��v���#�`��lmG��ȡ����^��u��?�9�]��XڇϺ��3Q.*ĵ&�,ż���:~�1]i�AM4@����H������v����2��;$Ꚋ��촷ogo0x �m����a�@��0c46ُ�_�C������B׍d�nC��M�wsIt��ٺj3}�M�a���Y�����{�6�,�Ȋ�gOL�!��1'�a�l-�9W5t�=����5���P�f�O���u˄߫������k�ҳP'��9+X�y�M��)��@��*���l}��{2�� �!𚚄;%��"�"�I�аx�K\k�`�����9]��Y`��xl'�p����>y���(���ጝ����Sڢ@vgMw��S;��{ݾ-.�	�� �\�����D�b�����6�����~�mZ[f{����#�%D�Qi֭���?}�?�Y��P�	G�<m�7K��Ad�ǆx�PW��T0A���h��P^
���/�b����_.}V�C�j�����-�*t�F_�G5���B�<�p�R��zN`�Ġ��ϼ��Q(�G������X�]���{�6䈝^a>��Aw�)�j��SL�;����U?��d3���z� >�.)�
�8��gp-��g0N�:����)u�Y��yFN�|/��9l�dC;���t����=pb��2�D��"`F@%df�����uhi=ў�Ϧ���@2O�=�q�6�K�(���{�������|ɽ��<�Y��j�-ķ+iu����@��i,b�J��#ys�X��gw���H�rɧb������
��v.�k>���Ν9r���e�U�D;��k���g\�/�2Y@֦@�E̤���t��BCV�/7sX����Ut6$����yG���5Ӆ;��Q������qH�v8f+�S�����)N��K��c>���l"?~�o�?���{/Ab�ݬ��bO\+�T��f�b�h���d-N�����}�.������������__�����k�&RF�	�L2`�w�f��}VN����W�~�i�L�q�C�tut<%���@.�L�����m/g���m#Q
�^S+���a��즡E+�i��������OϪ�=)��p�&�#L��W,�<YKJ�=���_��V���'��ژ�Q�~ɇ�������Ϸ2��$�H��8������ `a�V�,�M�r�J�k}�H�W�1�El���+�1K�5V�pa�����Ao��R����p;'�,ړ���g��@�:�{8��9�n�2��z|0�����(��d�DEY�C�-�.¼K������.�a�i�f����3�W[���N�����ܔ�`ç'.c=w����)|E>I��-r�6C�@Jʡ0~�a�6��-�����Q)�Iɽk.ߜ��E�3ρ��a�}�j/(��CF�K��o��r�
��*4��\F��q!cG �q\|���O�p��]��?Ɔ,5L��d'�,�rn�����|k� �fk�� ik�O��b<M��oS|��>�رwS���i
.��u\|�u�mV��(�+pd3�������6��K�j�_�d{&�Yp�&����΃[�olNw�a�<���f?�v{ج�ɔi6���qў�5���U�~/�����f�.v:=g:�'J�;���tԑ ���g,-��f��i4Z\�l���L��]�����Z���oy�K��
L�i9&�Ŗ�Rډi���.�!x��^>Zt{������\FeU��y翌��ۿ���oS�}��� ���V)Z�X�]���ܔ�m:M����fD����r�iΒ,�Gt�4��ǐK����r�s.Rt�m�X�N���;��CQ��zB�1����P������ND{&^t�D]��9�oX��>PgAǰV�1aB�v����������3����x�f���J�DJ�g��9���1]266f��.%�m$�7�E�Q�MåP�� ��ӿ`������	I�%\�6f�h��x)�ZK��H���W�#4yr������Ct�b�C�%��10����$w� Y�%(��ə��9����/d�4���NYW�����Ju�u��1���\?
v��4 cI���Q����{l��3�Y�,J4ў~�x,E)E�hU�x�#���"�[�9f0֠��"�R]��`�[�Uc�fl;Qf�8�qQ�-��I���h2g�_�ԯ�
(�O�����!s�#��0!9@��,�ȜRJ����+o3"`��/C���?B��x��>/�o�O��$�)i����/#Sge8�uW������t�=́�Id��[�&��\w�4\KY
kYVm�a�wa(�4�J$�7��Ƥ�ٷiii#�����.��F��$��2�g�GL� |i��j�d�S ���[�s��S�B�J)��$y�7��ucfU�g~�%�^�̂���
����^;��!�7��,�%i�}X���.ů�����-Xt1[RFG����4�����C���KZ1�F��VH��gff�۰�l��5D�# �+�ITl&��ؑ���^��m�/�CƦa�eo���"�Θ�`�);k�ӧݰJ��ڲHe�}�,�)Q ��ֺ��@��"�Z@D�@4k�����q��c[U��a��#��pw(�����4�|���+]E�(���q<�������	�\/�Xw����ᇶI�Rp��@
��>t��EZ��Hk�o�懐\6:4Yf,�0�O9r(��Nݑ��|�wh�C�j{Fr��6����/u�>��"ND��&#�ã	�C9�f�E;�f�jS��:��� }�������C�Q}H�k?�]���ѓ��B(هh�g�ډى����W0 ��bu��_M����-�nK�D�v�^X�VwB]l2D��YVp2d���	�S�	i��Y>�s9E�4�>,�M� �s@��k�z�&�3�&�%�	����&jsZݗ�+�aX[KH����T����EMb�Ђ�k���BQd�Ï�U)�MEv��Ԕ[�i�eO��J��+�-"�µ�I�e���s{������}=_��y��8��y.��RC��K�ݯ��ܹ~�_d�;m��9�'xg)������Sw�����i3O��>Ӏ��dX<c?�� ���,n}�����F_�1ڱ������1�,j����O������ĭ����Zȟ�� `�Wb��7 @L*�+Zb���4����Ԃ��q]7� <�?~Ïk�{s�MEI�/��1eOB�ƫ���c�\�[w�
񚰮YINM�uq����ڱ��$�ؼp��Ɨ���}��T�SǟN��iM��m���'D�������~�4_\>��USU�4���H�U��(8���%\�X	̚Y�X9��,� F��,5A/��on�l~%�z;�2�j����p����y��\�<)�w����|p��X�g�c����{� Uڸ����/=��M<�"D2���7��Ԁ��H ����: �;�]L��:�g)"�]�U7��B6!�c2LU㪳!�t�8Bw���%A;w�� W�3��O�`�+S�p� �����7	�	m_��.n�$��kݥ�6l���t]H*���L�a��
�x���"��XS�;|E��}���8%l�9[��hFaz��9F1.�Yyq���\UX���a*y�K���IcR펍���|��a�2����cC�ƶKr�f�!��1;�=�TE�b��N�B��yY\�o�j;(4Cq���ٲ
%I��&�����u ^�G�(�:�ښ!��1n
T�$�a�#.�a�SBB�p7n��%��{�j�K����?�6W�����ڲ��!���&J����I��tQ��'S��B�X#?w@�+k�z���BF��e[�M���M�E۞V�ꕵ�苩7��4�����Ma��q�`�����h�M�5"��9*��Fǯ�eeM��i#��
�^�80�0��`��N�����YQ�T����wBǊ��57"`��+*|}�S�(n ��t��Ь���5g2������&\�h�S�ri�"�\<��8��3�ρ��*4K��N���ySq�,��Ω������jV��>�р�
�A�9T�sϘ����� rp�+��0S�Ԗ�66F��E���=@�j1�e����	9��3��;   z�/wi��Ϳ���˃���0䝳���A���n���It ���5����Q4���Xu��E,�5��'�' �ZƏ�����}M�{�B�dP;�+r��w��Į�Z�a����f ���Zդ^��!����ᩓ5�����~�_�CKr��f;u6-~�����Rx�)<6��eq�:��ؽZ���#�]�L�М~�B�o9\K7�cՄ���;�����{���#_��q�O]�X�����-8�IղKLJe2�tara�"i�ם�f$��88�\h2�*�3��l�D�����m�[�\�I��7a_��y��9~=`�x�}�4:UZ@y	�
�\�q���V��KgXS����N�H����+�̨`�з��;0�~�755��wǽ����D�'�5���?�%s��O:G�AΊ}e��y���K~sA���1�Jw�Ahf*N�d3"-g?�r�?#��@p|=���4��(�c��B������,���Z~:s���&��ZgS���ťծ�p��߼ySa�
hH�ѐ&I�׫m�O� |�.�7���
cȯ.��p��[�]���
9@�[:#+��O�m�Cx��M�,��:
(J3h}�@��G�'������"�������)o0��m��� �Ơ"�iގ8��QD�$�C�l"��}h��dxj+c,�Z��&@\�|���1[f���d�y_�����P�K�u���6o��WT�v�{�]�������'�(��:�(2���E�� a��߷b=z��c��B��r�&QZ��름k�~hRrt��Zl/\D[�}�ɶ?Ο�[E+ڿ���I�5�g,U/���V��+R.p������K��|=�|(���%P撟�k!٤�yc���������������O\�Ӻ���b)�2N��t�H��pw+�Z�y��;GW�qp�*qa�W�z'�SrGvC��V[h�� �K�'��tuu��K_A"g�+&��?D~���3���טli3d����b6"zO�t)I��j�?4��6qJ�a��h��}k��V�u�������`P��黬!os��mO�#B\QzzG�"~�F����󙌫��<����C�Z�������H�">
�
^�lw.r/n���� �=��$ڟ�^�_
(,!����Ƽv`'WXF�9�����W��Ĝ��6(���_��u�$_ݵ�4\ס~�-�/1Ʊ�A�{ᑋY��Հ1��S�O��QS�A*��*�_ &8����n�
z	��B�hDhv�Yy�=}��rh�a�O�R��ttå�B��~$3��1qq�u�E8my?⸨���Im^���`�n'�@�촁�+�-6FQ��H}wO�3���t��b=�;t��ߝ ����:�v�v���Ut!v!���&�;cB�b�����5����������W^
�| FQ#A�YF+L�"�_@�h��$��j �<�W�{zyO��}}�7����JqW��8@�+�/�.��a��c���w;*2T[ʹ���u�=e��s���G����$v�`���s���A�ޮ
�sF��r"�*\TlR�<FY��|%�D`�����z�	xЛ0��d��X� �G�C�>e��}�� ��_��[xT�j�h)S� � 
Yl�/��rJSS����]�6]{Hdֲ=�5 *Q�!�p�q�6�m��o'2y���q���|Uە��꾝�ksN�0��n����صGNn��k�+�9�P˟`��3�V�i.؅�l��m�+g2p�k�O�BD�)��xp�8j]bNYO�������khh؝!�R,�BVQU5w;i����G�4�`�W�]�[�\��vyD�P�.�ͽ1�8֥��j��_&����|Ԁ�M�%p���{����Ԓٌ�l��`��/�)EҷM?g/������L~8�)I�Pm0)����b�3�ϧ�=��K��2CCh�)f�a��')2�MARQB.��w�ͬ��`]g���6��-3�Op�y�U9���Ou�}��L�5�[j�-���!E����"%��p�#�����Xvj"�;?��[�ȼ�+GpA����}��>+��5F�r�r����Td��e�;�ՠ�
��F��e{~�6һ�DPRw�jɄ���ԅ,�O�!h��(�5�n�C*.I8yg*8w��m��=0���T� �!j�@G��*��	V�C��ܪ���t���۔�N��H�
nܸ#�SFz�Y\�z��	ͤ�곴�%r�! �[╕�j׷����.*�z޾ p�9��ggM���<��n��ҢX�	j��.?����}�1��=���HNN��.�C[�x{�%[,�E�BW�N��:<��4�z��`aI��b�%�dP����:nf2{�Z�a婿[h��H[�� Z?�C��{��m
��Ox&��p��&�`�Bʅ �[vY�����Y��Z������=�\�&DL�E�t��.�q5�7��/���A~�ߡ;U@��(o�"@�,�ﴛ3(7��b$^��Xv��0z��|9H�˞�����aa���_�m>���&�0������]z��WɌ0��J�k g5I�M��Hm��[�鍐.�s* �ˈ�_%4�.H�,�K�C��H&��@M��;�	y�=[oҩ���'_�.K5��ג*d2���>��ٱ����L��#͑��D�丠�v�^"m\$H����ԉM�	�-:�@��|I�Kl�=�sir��0|�C��/j��AW�R��΅Ƞ;����8�=��t�D���g���l�Tܿđ\p"S�{�,.?�C����[�E��]M��NstL���o �VS�]R����1W�V��f��7���(�a��ꒋx���}��m�Uo� ?У��ǜ�1:>~��y�l:���<����:B�6VVVr
�a��S,da��e�Ux2���`�B@Ξ�g�?�	u�rh|���:o�vl��@��W�9�6�j(��BW�t���<xo%Ze��@v|Ι)���m�������rkH�Wy]~{���K��Wқ�}k�Z��S�T��t\Ѡ��p#i�J�_��ȹݽ��w��b\)"��M�g�P�^8��S�hK
(\��cɁ{GRw��\z��=���!�c��������n��b��2��8��6%��H�,:5���H[��-��1��U+����@-�8�;�ї��wR�������X�X�~�4
�<��\w��Ţ�`����zcV[i{���*\oӳg�.k/&��0��Z���q�]��=��g��yά�灓zc�o�\'+O<�l�J\��%�ң��<J?�Kd\��n|
�Ӫk� ��</�_�����!B�����wkD�+w��ʑ��Ǉ�X��S�g���}3L�D�ThJ��S�#��,�d���a��+�H��M
U1�:5��+7 ܙ����g����y :���X�p@U�R�L�_�]ۮ�3���6+� :�0+�Ӱ�]�;�3��&a��5Y�9�i��ͭ��������1|�7o޼�+y�E�ݨ\m����wa���;�����~�xZ����G[ɢwi�Ϥr�K�̮#��6*s9�!E���`��9�ӽ�j�T��M���H�"���Աy	�BD�p�e�;̶CD��q� j�z�XZ��>��G��q���}x:.�����Z�e�_�$.��o�Iu��ڝC�:��8����´w� a3�)W�o p[k3�l��]�&p:�2�i"�`�#���._ %��$�}G��$9�q�wAy���u��T�2���>|�DKCp�U�{��5�f��KO�ڈ�
����Hc�`}�;�ru<ޣ�g��v�;$$�7{ y$��A*�ޥcq|��uPR�l��=q�С%��,��pz'F�f6oI7l���G���*M^y#	����ŏN����/�9$�8�-���Z����5��G}�4=Ԭ�[�o�qo���f �-C�?/tI������q�����|<2�ǔ«!N,L/��x������cƖ��������,hb�d�?rUk@���^ rW�C��(c%1��V�*O���zx`��U�.��34o���M ��9` ���[t�vA��X�uy�"#��&��0z~� �&&&�1�=�� km�8�#`Dox���u�{C0U�Jð�Icu���Z�����v��[��92�~֔�x�F�[r�*q�,<��-��	Zz�r\;c��?|)A���-���t%F���r��W6~��W��D7���t�,�'�qǜM)}�u��)Y �z/P��v����\�.�@�u�MZ���9橞�d�r�~�ܤc+uϦU��	�������[IrC�������=����hw�\��_entj"J,!����U�Z�	��*�"K��4Q�4S����
�c�W�
���A	�/-"�!��"1�i]��5�\��h�ϻ�mC�뚥�e�q�mlZ�QZ�5U����Ss¶�����O_ ��]Z���ݩy�5�(�x+DN�#!X�ƪ��7]�^�����W/�J��+2��-6���˷whh����*�#���z��+�B$���;`̱�%R� ӑ'B�bmN㼞�����ih�˺��<�fP4�����M�;��
���A�?���f�%�D��#�"�����	�3 Lԙk��K������Ca��a��;i?�Z�$[�EdT�w�{���C���Sj?�.�j ��fB�����	���Q]mM��k���eaM���]@?�9;��q,�����R�= �u�#\eIO��7fgu �+��FЎ�?>�ϲ���NOK-�ҵg:t�o#�a���d�f�};�<^)��'i��Zn�!cma7��n&���KC������U�{փ�oxΠ��H�|�U�]zwO6��]�����%��s\��z�J���۳��0xď���	�����ަ=�RC��@.�Y�ibb2�=Dg�;� |����Z�5Li*��ڔ��I��֯&�Sn�8cC�eh����c���Kᙤ�f�ɒ���?�����&���K���C���`@^��*<�4d5�!��L��ܢ[�Kj�s:w��W�ܝɇ56����������ռ��"9�r�$s^��s����f�~j�q����
	��4���0+���b�-4]�����/��$v�J>oY�!��@��e{�C�q�p�������g���)���Zڒ[n�E6���L��_�5M�u<6xc*Ʒ6�g����:�58--0-�Ub��^š�R7��"�㌗��G����Ɩ��i����K��.͹�x
SM��C�I4X�g�)��ɬ��7nv宒w)���L�6X-믎��IvD�,/�5Dw���TR�k�yD�ʘ�O5��픷k����Z�0dw�4��8*wFe��.#��o���Bu�L������RI�2y����{��Vk�P�6�����0~���_^v�IT�v�3���Ů�7��<ؼv:r�#�g��b���q�N0�3����#��f�z�syv�y'�h+<�,�SG,����/�tq�����˵�fU�<ciU����0�+ �|������,#-��;���9r�t��#��*@Шn*q���
���zĈ�=rK�(��V�+�(/�����v%g �����7y/Z�����M���r�.�G~Nڱxx�����E?&s��_��z9w�r��@�Kh#>>&�D���M"1�X�n�^���h�A"���pQapo# ��} �vu(V�k���wv
����O*5CXgX�����w�I�j^�5(�"6\tq�`2��o�/]駌��rj���$��w�ET�Q��u����ٱ^Uٞ h��&��7]N
���x�����0�-�+9��,շ��f���`��Ku�b��"_`v������1�
3�? �e��@���8B��P8��(EB^�-+��#:x�:ٞ0�}`��oU�ǉsVC���۪++����>L.,Ց������f|h��;���Ju��LJ�p;طN1��d��Ln��Ƶ_�v�c��@<���11�p�7Xݑ���_�Å��׉6���$o�mK����o0��XR�Wq�;��umY�x�%���L�9�����X��r�A-��|}i&
{�P~Jh%�z8�!�q���!����D׶�c�^k�mi� v6TV�B�����cX�'</�t�y��\w�mu�"2��2~I�r����� ���C8�J^��1�p�2t�Q;qMS �|��u�:$:�3���pSY,u�܋�>��L�i֣ȝ	jj���9�C,��_BBB��v���K��'��{�v������J4t7�ӟ��{��)b��)��#�� E��[�t�`�ՋՄ�.[VJTн��"D������S��?�n��ƣw�C���/��X��J�T�t�[�d���l�� і��^+ypƋ����s�AC����=l^|*��P؝�l����F�LF  �Z�)n�"<y�3�ۂx޺��zB�ڣgjb��sF��I��~��徱f���-����m��I�f�KS���Q�yt����:�Y��Đ����_�S�J/�������жO~�m�D���,�;�L��U��9�D���8�Gi���G�$b�w��#[��65��4�Yex�"������lI����
3��(������+9%�v��
��Uon�1{a�M�'3z�쒷u��'Ak�i<��c��Ќ���>(�!����:��ǟ���(z�*xa||���4�g���\�����:D<v�$��:����PF�(d�
�����&�u��U���ӵ�5{����[l�o�ĵ�le�i������9�M��y����g�ɟܓ��sIwQ�t��4� H��Xj^/a��f�A>��z��V{qhyia����{�Ɋ��P�栰���ٮ�U\®����a	��~��d����'��R�υG�m۶@�� o[��	<�)�6p^)&�/�8i��Ka�!�Z3��$�O2�Ļ`O0*

�p��:�����\��,m�G�yn��y6�3����Ej����-Iy�%��#�pFϥ��03�b˚څȢR.�b�=C���^����
2��D�.�m+������
�n*R�����
�b.�uu�����%�p�X���3�������`CS{ǋ{�6���~1��ӱ�b�r�Z��$���^�1�����b�J4�S�&� �h�*����SI�'�מI-��U5�,c�߹�mר �����P'�8�Gq<A����m0��1ƭ!&c&4r���(�ͧ�C�qX���(������!�����ab�h
����xd�*�3����d�`q��}���b38�$}�&�L[w䅩*�}�0�.�3�'�*�_�b�b���c��7b��9��H��}���^h�@�a�2Ĥռ�Q��I'!�d�N�{�K�/��2�"}�U�D-W�N<�{J��O�=Eyܡ���<eB�uhI�mA�0y�:����ߛ[�V��|�@+s��z��[��"j�"rD�p��e�/����ix��+�-����	����)}{q�?� OSST�1���0�4�'����\l��R��Jg�z��j"�0��˵��B�c���f:�Z�8]Q��\M�왝]ߪU@�6��(.�OVWS%��S��Qg��J��?�m�ݚ�f�/ҟW�=�罌��=l����:X�����ve���j�!2���|�&n��C�i��3 �#�w�:p�?����(.�p9&r���=J��	���2�������m	�0!��˱���{�2!��C���+G��(�e��M��N����N	�7?�h�s<gY[���F�80�&�B�;��~Z=$=GAY#�î_��/#J�R��o��[�,��+�u�]m/q�c
���%ݶ{��s"���ډ�Վ����]<Vi�SU�o/ �U����q�ni"��*��ǌ�j�Ζ�o>�Ù�E-�����v�����/_���8�s���+��? (AۮG��&|d�$�H&'KP�L�G�1ׅS�Ґ@%���b���P���:3Y:Q���`jf��>(��Y�Ϛ:�%)��

��B?!�)��[ �)��k�!T�^{���i,z��7�1�����*�X��v��.�a�:��==�:��튣�3CM�K�6ѭ7��ѕ���c���[:=6t^ii,�V �\F/`P����]�q�v�A�8�Omy�ޟ*���g�n�r{{{��2D��;wdR�-��G3M~�[��I��ן0R�xH��^����,z�}Wo�Y�X4�h�o�4]�W�x�3��d�xP-����z�c������*~�X���0L\9���d���q�Մ�K��`U�̍!୭����Hc/q��B�(��8�Wr�������������D�1����hǃo����H�L�t�l�a��G`5��ngˬ���-@a벦�R����������j��$�k���w߾�Cd��x�Ӻ�C�����h��G(}��ޝ��R����:� P��v�B���v��)}�q����ݾ��zy�����%��j�u���9>c/��J}vS���G���{�dr�Ԁ���x��M�BZ-���V�J�/���jB^��ʁd�ŴD�^�b^�I�����j��g�RB3�s=�5�#�fya%����aR��M���\�&-��������?�<r�R?!(t�Bw�#uO�Y���K� M���&�Ů1�fVS޳,�J����ޖ� ����8`fN�=�� : -׆n�/ �y���?��(�(���_���{t� ��;�^�b�<	�x��!�$��,��TF�튧��������B� �^��Ԝ�;3����� �!�d��2ģ��㪼�"�?�H��}x}]d�Gy��Y�I��\m�H�@a�u娈�u6�|bf����M�n[�x�#�҂�!�I�6נ�9 �0�n�,!�yJ�\5�N��`E�0��WL��ů�G@4��F���k��E��̿j�VaGH6�7�b_.^P���k�w�<�n���{h��o4�%%�r��ʑ��%D�sV��2�8�X�!Z���IP'�n�+C�Hs�e���"X+=��S�� d0�M%����7����[H�����H�;Q��3V��������]���~az�,�0y^.;���F+?�r�i���i�|��\��Y;�P�H���-/�R��@�z0&zsZx������|�n5�20|.�����ʗ����TM�����_Z��z�A7iK���{�6���ߴ�#B�ȼ��m�_�rō$��U&?�M��	��֖t�|��R>D�=��u8��4��>Ы��6��I�Wӂ:��/���o��qx�_�Vh�\�V!�L�yU��K�$9��
�5��_��q���B_�Z������[3$�?~��$/_���Ro��Й��I���.���������)��Fȯu�+�=Z�7�C��*s�~wh�ވc�,rcFF��-:V��ϰ���>O�~ᩔ��a:��5zz� ��/�]OY��z3�h˒���㏑��_Ss��	!B�S�s�-ܩOU���o������5�=���{������N��|�O-�������
l E����
(Nj��~���6cc��=L����43=ʱu�֍B(�?�π�'�Lz@V8c�^8�/_m�������5A> ��g}�Ȳ�
�j��eE85��aM��=�Q��݀���� ����-�4�H׻��|,B����m$�o�H��)�s%��G��U�� �+�kJ���:褷3�矿��Q�Ǒ?~x��:����)}.�c牋nxp���N�@�ͨh�a�o�Tÿx,�7�>���7��� ěo˵��E�/���Evvv���=�^�JއE��!`��|k'�X� v�%jA���S���P�AC��3�e��x�Y���d�Bj�o�N����;e����T���r�������V�Ic�`/�d����ݖ��P�.���)~�]W\^��ۆWq�a����ĉ��c�C��9�n�-H���Tg\�Uޠ;n+<�_8V�ጋ�g ��_0���?�dvV��[�@R6.��z(�*�x�u��2�`����_ӆZ��o���;�J�gb�A�*����y�w�gu��n�}�.s����[��T�.�җm�Ջm�/f�'�ʑ�D#������>DD
.��X�K*�H��g�b��bl��1#I���R�0S�O\^s�eH�~SSSƸc^��^��8W�Ԅq�y'E$o�Hi;�/J�y}}H-O�d���Y����8JuIls��� �f������������}#���E��6�����D�����K������2V�dj����{~�>���_(�kJsraiE�rkeu�O����%��L%�:�H�5�j �O�y�������ru���q���p�.I��I5ndl,ѣ8���0�ή�f5D~G�x��6\,��3�ƏXk5q�m���an|qS��z;�2V�è�u�c�D�)�Ü����8�:K��[!?vg� ����\�ę�P3X������@�q��<�˨=^ ��I�;ɔZ��W=�⮆v�ƚ���{M9�O�~ ����N�x�.���$Dp�A:��#1[=���8����Y̾O���
�\I`�g�D_@�WLb��8����/�&WK[{���46��Џ�]^tz'P��L�K�]�T�C�W�3M	Z��;؂�&?�����4���+\������r^ԟ̛�tY\R^ �"��d|w������ơ�{_F5iuz���E���'�\�n2�8�"������ �b��<�\/�����j=�a=��XLb�^d�-fs}ƺ��$�a}z���Q�[ǟ�V�jx�E$�s[�Bd;�����I�REւ����d�������� �ݺ:vN[�oo�Pd���)�������XP�u��ˌ����D���7�����|��öm�d� -vB4K�d�X�����w%�7_�vK��|��Wg.JV��K�r�0�,..J �K<�j�JIި��>񓓁�"t�/�UD�ڢ�4�q���N�tU ��t��}�O2*��#b�8A'�� ��g�poWw���~%�@��k$�B�ڣVu+�{}|�!N���{a}����������ܚf�d����K���z{���#�S�^/��.�	r���Q����?H�� 
�
k�4+V��]��R�]!k�w��������>�n�x���
��R�q����^��L������[���F���c]Y�H���͗#�#��� 9@=W�K-����?�J���:c� �햞��K��4�����li��q��D�̸�f�C�ALTԘ��s`�G�#`BF��;���{ʼ�{�+ ���]�1l�����А�m��B⻂Or��$���k�ׄ��jP�Z;$�*��������c�Tg�7�-8�{RqT�ƕ�����u���忓i�߮��BV݀$G(挞��ZP逨�-��g ��ݺg_����l2N���i�u_�T��$)f���d��ꙿ	B�R�#����^��C����Kc�_6�7Or�>�O��F�iꇄ�C�Õ�ǗS�ňDVÕ����f�	���V�\���"��L9�)�s�2d��Ц{����ԛD��~�x�|���"�n�*o ��y�GS|���w�X@��͇��vNr�7����It��8��z��U����7�u��ߡ��4}�h���ć$��������m2dҒ4�{�F��3��i�����^��WU"��(w�f�{i�D��a%�;�>��i������5��H�!�+������R J>��uq�_W!$���}�/�G���H�g�����bN��@��-��`�S��4_E6;|�(Ib\=����g�'O� y#��,O��ΑH���� z_feM;�{p�����={���0Wr�7<��A���᯸�����Ĝ�U���DU㪧����pE���Sw�Cpsr8}��(.�s�d����p�n��M��c����7)��C%�.t��{ā�p�S���G��6�)���A?*
W^���,Ǖ�����J���!�yB^����V
���;K���2|���	���>=�k��t�W���C�:�y�H[p�9�7?���=�T%�m�����2�u�K޵W;H��*���d�����[\+�Y����p��Ntv���HL�CC��Oh���_�L3�]6qq��&��ؘ���Rv�-�$9X5휧S���I �J�(O���"�Ms��ϲ��NLL�B�ny�3!�nSn����?��Y�[����� ҆�f��:�:Vc3vK���y"��=]���������x/-#V�;B~�J\����f�%AA"���A�dO�89���X'͑Qq���{�2B ��o>ѦK���YE� ��P	��ςX��E`��׳վ�\������{Z���
�WPs��!q��ﭓ�F��g�tT��q�8��塗�L��02ח��)I����P���TˬO��V�5m�]:ӕ�.�$=�?W^�B�ki!_�(�jJ�5��N]���8w�IbŊ�:0�ZDƯ�Q3s�ڂ���>z��+ql�̰QH�wVQ1����h	%��}ՎZN�����k}��2.K�Y.��k�\� L+�~WI����Yᇳ�v����u���Z��E��A���|9v�>�3��HM�KY7B�Q�����)�UjBg7}7�d�g�OC�7y>�hd�t����l��+���1^�u~S����{Sr���t�*ڹ�����-q���-D$�	��9?�Gx���\���tmIIɮ�۪��g����n������f�e-;S�{j���1[~¦j�ňЎ� �fgm'B�Ta��#�GLT�5{4߀�k�1��2_�x���lpA5�-7E��*!�5���΀��U?��ʉ�nl~2k48L�9[�N�emgM4���æ�B�>!��٢Qv�i���k����Z�-�a�tC:���@;/�C�6�"�V�5�)}sc�L}5t��G��I�������
KW�	˗#O{�N;k���S��>B/��#)�&cUyGSSSCl�;boo{�N�?C}$��H+�4�m�7�n9L�-yYÚ-1�f�5�R+���mA��=
M8�.�_e���V���N�-��{%Bo�Z���������v��`P���w��^���K=�9���6k�h\^4�>֖5��w�?;�סSb�O��o7��l!���,���J�?��Z�[��jJy�W�ݧ�l:�����x'��B���b5��b�Ē�k����A]�y�
�w�qL�N�c���(A$��}��1���hG�6�W]�z�����9J_��7q�jBޜ�@$���@h�ټm�7)�	��z:��ڔ4�q
�šU�*8\{��o��0mr�9�(ڃ���,�x7UCV�{�� 6L4ڂ�pa�ٻ����ރ�P�.�8�1�?p�\`�*��a��s���"�G�kfjۍ�e4�ߢ�;o���.�̷�^p���9���`m�w��\���|�=f�ēi�޻nE�|�G���7�?��hA���u咠���	$U�$Yݰ��$h] �e(��QNe��l ���rq��3g�>-8N&n�i,̌T#��|����1�ݘ��8���_��C� |\	�4��M�������:�X�4dܚ5�����s8��LksP�tlM���wĉ���s7�_��<�1Ϲ"Fp���xM����k)�FXe4Л��	�5��{�-_���d��ҡC��"d���8�OEaJ�27Z�<�[�I	����G�0#��oj�\��$��LOmj���v ���EL蠉V �1ڀf֬vӲH�/@����U&g�>�����So�-r_7<�P���CZV�1U`^��O��ǬL�(�.�Ro?]%H��-K:�2�/��|R-�1���<d2��v��9C@�M�>W��"��$t�M^ֆ�kE'�]�������?*Mj\���`l���(*	~l9�����gC����N"��9��jy#v���W�P�DԆ]��p�����>_��;�����$��K�	?��I�;���M��� i��=[N��])Q�� D�)o_m�=V��	HV	LJ�A�F��(-:j��__�����>�s� 3��5�Q���A�o���O�nL���Y�p��cq~�4�-�+M��}�_�Um���ܤ0!�p�HW��B]�� !\^R7~�,t��	g�y��A|�5�[��6K���dz�S��WT+n	9h��;��!�s���M{t(}�c=G�|GBx��n�h#L��J��y���|�����_������R'a��Dr����������u%Z������g��D�9*��>����0jfg*��0���:��D�J�~\�,و8���P> ��_���J�V20����+�|/�^{��9��W�����H�U+��`
�#��X��y���(�	&��Y��Y���X�Ѧ��FZ�]ǥh[�z�	��㽰�gP��@�u������?idE���L�l?=2�\� ���Kl�9�y�bo�Y�D�Dӕǩ�������X{�UG$ژ�'|6S��T�[��<+n�nS[�C�О�ґ�
t�4������k��ٝ����%�mi�?��A˫%�ꮩ��f�Ʒ6~J��5��0B���r9�S�B"A��J�eV�P˕06J�7���V�C/dO*�coq]�)�?`�?0�m���vN�sB�{�k���{5Bt��M������v��joo��AZIA�"���j��7��)� 4������QvQ���Y��=)���?Tݸ<�z���(�� ���(˟��m��� $U��s�"*� �ݪ�}	�X�$hJ�����+�'$�������vA�(;'�;��%���5z|�Y����^���nP症0�;�����B�k��_�_�L�./�ޒ�3�~��0�n���H(�r�#}.z V� FL�,�i�7�U�5W�hu��Ͻ��Rn��r��՞�ű���w��=�,L�����ڀ�J��_/u��h����8*x��9SӅv��q�@��0��_�kl,����<N(2�Wc�^x��M��Ν-->v+�iW��R�pr���Pe�B�3u�i�&��D4�f;W�	��Q����aK��&�3����Y���ꕂ/�U.#�m�z���K��u�\�ѭf�tq� v^��̀_�صN?[8=�,�p�-D� TQ�6��q�����h/a0r:�o���K:=��wޢ�@�Zbg��È�)5�o��B
L�)��O�/�sQq�۸i�Z��8%g�	�ȩ��nyY���B|g�}�ݷ�Z-4i�=��Q�$0h���ұ�h�@��Dr�۪����VWY)(m�8.�>a����{W�{\?S�"Y�`�*C���QQN�j��憒��V7�a;�A��H���,�wfm\7�e�܈c/�7��7緬���@F���\=�Rc٪t�NH�z�dk�Y�L�""�V�k�6{*�.o+��b���x�Ҹt�:���q% 膗�.��C;��i^�8	�w��GK&� Z}|F/���h3���x���k��ѕ�m�du�!���/%⸩�|�*B���(}��7�
���c���:�7�~ӣ#d��d@$=�Hr�p��Ϣ�T.&�l	 .p����Z]a/G�"}�}�H\=���I�V�A���[vl!u���=��cQ� /n&a̶��!N^h ���2b�'��@z!�٩u��N����Hj(o!��|�@p�\�Y*:�w�s�ه�r�O5�e���Bd��֠�l� ��"��a�Mt?x�N�A�
ӎ�~R���ԑ����dK~J5fksK��3��˯ �+V�`�����S�����ϴgo"�)U���Y*�koQ���#!�$��F�O��ᓟ�\~�����ĺ����.%��%Y�O�5N`��0��r(�ң�:�&���'���y!��̠jP�1ݗW�@�B��}�Î�8N���!�_Ȑ���Y��fЗ#)�D"�I�w�O�+�P�p���F$h-�3�����O~~o-ۓ
y*��︯k�' f�������;�*���ի�k��Tm|D;_0zn�kY���d�ɬg�X)���.�=��|�K��)6�nN��֨[��U܏�nDKF���V������<��LIL���~��~-�UK�p�+���5r��F���m�?��r���>��	>[�|H-��M���[��Tw�[9����_���c���]bnY99ޏ�+^��:��+� �	^�yx]�9Lg�s+��>i蚏��ރ��M/��kõ�m��v�P���|���%S���O�8���� ��tyOKIs/����5���'"5������A�8>�'�"c��y���Hcu��6]'�&*����-�}/8=���~��=�a��G>�!���x��+��p1\=K�,vZLH�
˵i�ʙ'U!W4(��wRpP%�A]uֈ﬏U�	k�3Ȧ��G��L�Χ��oAt�TH��}�-��}�k�jt�æ������BDdP��ƶ`8���V	Ll0|٬pc)��0@t�h6� 8׽G��#mJ|{Vf���r�o�J�OB*v�<|t-(+`��0�aY�W�=�-����4����Roo��X'�AZ?j���m�2�M�J��h�m|��3Я7�8���(q�YH����]У|7µ<ΥR�-�~n�[[k<V��^�^�n�d�<��M�=��� �5�l�G'��üp0���ؐ�f�U��Y���R�=�U�Y�R�K��Xu�����b��Ǜ1���T�\}�����g�t�9rO!�#��O�Hw������Gq< �o�B� �������L�Ma��*��ϥVE��l�U�#���Q?��Ԓy$�����Yy=�S�	�kS������ޒ1�f,�R���a�S�}�~Z��A�F��O #� "���
g�V�`J�_�sBv�m�pVk��DZN�ɑ�sb�G��j�_ꓞ��ў�]Z���Hη��!��%eA�����!�Ç:c���2�u#\�Y'PpҘ��=r0��������;��.�z[lK�i�bL<P�5+�H�7W��gTU�)J~"$�6��L��p~v�~�mD�FDI���ް~�^�m��� ͱ|����T�U��QJb���Y@��tް��)�;CQ ^�k<��w��Q*���!'�%��;�"$����Βۛku[�����\�#.n�dɪ�'(ّ� �yp�}��Q0����A)n���O����I�`7' ^���>S �~�qj;�~Nb�\�?��&��S,,���M6��[�KSQ��23�2�jD_��̙IEٴ"�)�Ԝ�"�,]YHXQ�oZ��t-Y-h��F_���@�U���Q1���}���[QA���=�s�=���9o��D,���v6�w�-4	���s�$��;�ޕ;&xdR�����ba0�lw�:X� �X06�ֲ�g��~-k���=�3�4��יć@�35�^�{2`�xU�� ����W(e$��!^N������OGg�)���Th��-e�A�������N��d{<c���2���mͽos����C*�	�����c}��J���a��b�W�V��~8�Ds��f���@3NݺX
�-+]��v�u���t4Lf�M�q�����+�ذ�a�_���������%T�����N�[�:3�A��p�3���)
Mk&ثA�����ъ���l\j�� &�J�s���UhG+��3x���Go�.7T9U��|:[�����`����DJ	Vg� t��5�ܣ�)E���KI��Qk���D�
�%��q+֠!���ؒ��z���������q�Z����̭s�5Ҫϙ&|Gøn3dE�d�򉼩j���lyzd�8�<�p����G����f߀|!~c�-L�_�-�	��0���Y��~V?���?gum�p��j��l��Ɂnb=�e2D�w�{�>"�Jm�.`'p `��]�1�3>��B��2e���C��
�[ <�(���[��&�yf[K=a ��)ĵ����XD�b����n�{�*/ivB^-o�p�znGx�n���(��� ����Jct�������J�<����pÖ� pPS�q����(�3�ʴ]��<� �4r�Q���+��9t�Q��Z*а(�ji��x
<��� �P[na����N��n��x�/Ù_�Y��mj_֡^�=L�"�:�=*-}0ѶE�A�5���v6d�@Q@�iE|x�:�b����G��jJ�&uF]����Â\m�h�#��n=�G�H­E53E�Xk"lN	M��_�n�;�ZD��9߾J�->�OX��w���e�yW����'�D�V-_�b��PK   �c7Y	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �c7Y�h�F  A  /   images/cb0ca54b-1964-4771-904a-f612fb73280a.pngA��PNG

   IHDR   d   �   �8�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l\�y�]ޗ(:���D�uR�]���ZM]'q�&��Z>MѸ��nݢ���h�(5Ңhc;��I��)Ԋ�;�uZ�e�A�(RI��!^����f�����ݷ�%�����������̛�.R�N�>-����|"���F�'?�Q�Q�P�J e������Y����Ν+R�R���f ���CY�R#l 
��栣(�d�䠔�T��P�Q���쓨���S�NY�
0�b�"	D�(KP
��Ԁ,�.U:A"e��6�W����;�υ-M)̄��!���r�R�La��!n�u)�E��G�e�Nu��f� a��~�e/�m�GY+l�C)���|$a��g:�WP.Cy�޾� %��R!�X��Ua��!�D"���;7==�ppp�J�7(lp��	�P2�D�e��m΄��T@����j�?����v��/;;�6++k1��j�p�B�9�4`(-��+�mg^Gi�'�����!��7����P�B~ p@\�����<���,����������v	
�`�8((��By���K&(I�F�ߊ�u"�TXz_cTLDЇ���QW��S�%	sQfARN���!hi�R��w���k��`�@I
 
�RF]X0�0������򾾾�J��q_`2|RQ$��?�/��f���~U֪���ɛ[�5�y}2@I8 #N�&, �,//o%�+HKK�����TH[˽������C�Q�B�9Ch%�{�\	`�AZ5o�@�o����q�Ii�3g�H%��-0���*a�'dLL�����9�R������Fn�D��^�BZ �\x^KQ�0*&��b���dwww柳A�K~�(]��sJ MMM֧�\�ޔ3�d�nڴi+�>��E7� @��P_'� ŧ�E=' -�_�e��KbІj�' �>))B�üٟ����`"UW� ��+�Y~��(���������`D�$(��:�٦4ؔ�s��m�}/��"W���H�$��36���?J�=I l,T��{ɟ�
۷�� �Tfff(0FOS2��� �-������`��@I������7@cIj� �t�*�&ı6� J��H0hDi;�D�Ҁ�a�&.��p�z)xu�ۼhA(Ð�Ϡ����. ލ���죇��!d;i{֡��!%����R:�
����-�)q�pF"��vآ#^������ǌ{4)u�t��e��H %�ˢ�\&�G�A��Z����d1j��h=F�P�6$�=T�hX7U�<L�ざ�1{�l��9 Z�ragnu��4z{�A��{dl�O ���!0N��H����M�)����r�v�3~b:U'	Ƒ+QJ�12��O+�-h��)����(3`?JEd0Ҡ��(��~N+�om�� ���<�8Q6��8U @ F��v&�N�� �����2zO L5pzTg:=�l&�Dd�*�h:Q�kb���j��-�N�d���TW ���l���po�&$v��}�3VC���-���c�AxV�rb*l ���f�#Km�Or���5�y�#��v0<��U�*�m�N�'��R�"1v��d2�G?�y'@�$�ľ��ūJ=R �X��Q�S* F��:�`؏sb����)�W���� ֗�<@RB�����>19�6Dx��z�������Q�j�'«,b2$�?�@��׀�"��P��'!y:�&|��F�Q:<�T��K��]$�� ������G�\��2�Fi��dP� ���Pτ�I�0hJCo�R!c���2MC�c�	0��w��ܹs�>,���˗�[TTt.�{�K�\%(<����͚։#���b_III�b`$"��������Pw�yԓQZZz�2u�����9s�����&��E~[ОN/���HT���YgϞ�&^�:.���z����7�p�OM����*������;�g�dnNN�������q=��f���C����RH�d҄ �tww��LɄqB��>|����� 62�t�۷�#T=`��]�v#%���Ou���Tv����ӄ ����ϥB!AЉ�<r�Ⱥ���c�����-�8q��<��+�k�׬Y�*�U'�R��n����h׮]롮���l����
�����疘#����������X���P\��+�JJ�����U�V�����UIA���ر�؋҉�j�Dܔ�X:P\�ۡ� ���~
	;�����ח�}��o��MJ�E�eECтH0�����ת���@%Y`Hg"c�֭�Am.H0H�
�h� .^���%K��\�f�AW`|jsq*�A�Ҁ,Z���+V�V`(7v˖-�ttt,K50HS�*؋M�W�ޮl��� _�W�:� M9@���!z{{���!�AzT۶m�bkk땩�M��)��ٳg7!
�@Կ����:����������SҔ�`̘1�F�A�5�cj����G��"�Ju0HS�Q\\�VSSc��"y،�S�N1%R����DQJ��,gB���pm�+Um0�R������X��p�ڦ���@B��6����333&�|0�Cpoi��p�|s�������n���P8<<�'/��&ـX�|�dF8�O�����j2�!G�O�!���!D���`P�>���Ո܋�j�>�*���#ZJ �_ �����`^V�s�PF���Ա�)Xǳ�֡���jD�"77���3sp��(�|�]|����J �� �<t�P�{Lb�kڞ����pFv������⥗^��w_\7L8 T��W�S'O��?,��]UVWPP��i|
������r���'%e�ƍ�{��~	�#�r.>�`�'bB2���6m�g���*�3�������ӧ��1�Dn>�\5tp���'�����Z���~��и	� 1@^~�eq���t�D��2�����{'9�F`K!��)�� w�À�}��v'�$�2��@��#\NI�/�[}�E��^��B}����*%�B00�
蝰�SD2tb�Ҡ�+`۵�x�߻)%��b��S@�;�(�{�d�[�6�n|	ݘǿA\����?��},{
Hvvv�5�z��!�6�a�9�"ˠ��u��W^yE�u�]QU�) EEE�����%�ħ��A<���ܗ����3�׃�ak���s�Ԉ��x*��Ə{���ȵ`QW� t� ~�c�S��;�ݬ@��]�������`!~�ɍ�s�C�Z�	�IM!�m&m�9�D)mg��A}=Ѷ�3@�2`v6DFtqqsNN��`U��r{
k�������p�

��nK-��]j�	ڕ�X���J���y�e��8��n�v�W[[{�}�ܠƗ̇dT�*++���'r��\�s��JrqG�X�Z�r��>6௮�N�w�[9;��?�ݗ7�f�D�ZE�w�	rcL� Q��3@`�Ekk+|Y�F��������=��Q�� �8��uww�#��]W�)�t�j�c_���,..�_Q��i �iН=S=R' `8gA������?%rY�R���(AHI�ta��k	���� ��%��\�pNC�ma������%j�J���7�|^2�F�1~�����|	'n�b�����KP T���+w��2��+�3އ��+��#��P�����w���:�NL1W���t��"�|�^6-:{�,Wd�1����ӧ��+`�4�Ch�BF����"� ��\���G!L����l�(ޅx�G�2כ/���p�677gp�u��f̰.e��,U"&���Ioii)I䫁"6 N�"ҲS�:�u���!��h�P� �/;��C!Eڒ�dS�����`�w���b9mkW�Ĺs�Z�W(G e�	��C�����)���-�����xYYY�+k�
�O��h)!��!\iB}ʆ���q��:TU�(� D�AG�����FK��p���%%%�)��ȕ�#_�4٤E�?��������[�pa@�G�l'��9�[�lY������Z>Jܳg��3v���+�.�:T_g���5��KOO�80�@���a����#q���6�F|޼y|gT�����������j1s�L���'�M���lc	��ɷ`/^��H0(8�'���ӽ�1��V��Q}=zTvl���V�8��QGP��SlE#7}���TQN��g$���P��s8��P�Z�*�x���a#KKK�r�������5���JUV�	w���yZ���}qD0��MqX,� 8�k��>-X� ���L
���!�>�G���*P���:�w�^��c�´4�����܉Ɵ;�Lc�M�^$iN>h�l�'��?�s�Μ9�O	vzRtH��<z��!!�7y؉�_��+W���M� d�Nv���.�@ 0���lV^^nƎC�1�Q��j�Imܔ��+U敽����ol`.j&�s9O&�����Q��ީ�N��`(�
;$r��X�U,+Mt�fԎ�,��!JԙF! �+����DG谟#T�s�q� &	-���rb:SU&Y��z��ĲzH���}0H8o_Ku鳉�ca�y_�LZ��S/�r<4J 8��B�z^K�/_�N.Rd���_�7J�dHMM�%��N�q����������3��t)/��u��VF�M#* �-}�b#U�M���7N3U��
tvv�.�	DEE���@�X?�Ƴ���J��X�"nz��-�Do���>����2��%K�9�#2@�ljjb�����f�� (d�Rj�˵�K���)|ǭj��)=A+x�4�  ����H�=0A�A��p��=���</O�� 
�N��ןm\�f�ZF�A���F���1J9���||�ɓ'-L���[ޙ
,y��A}���.MT{�^�S�Jq�:�������WI`�g��|�P����ӳf�=N��<UY���v��|���:�`0A{sJ2��5�L�����Ĭ MT)1��g��ըU.�ܓק�7���) �3�K�:7�z������	��G��=��hԾ���Y�ٹݻw[^�ڵk-�n�)���8.�P�%�HWF^3�]�0��|T��|��S3}&�;�cǎ���F���4~za3���>-&p�֦M�,�N�F3R�G�D�p$:S.\�$B�,�$1T���ie(��4�6�^RR6�$#�:c"��@���S�Ȯ��OR���؉��� ��&�9��;Y��$s'KZhP?��+��t��~Ω�ɶp:ٓ'D�A�8g`�D	%C��Mi<Dُp��a$�m۶�֭�s߾}�p�6�������^��5�F7ʧ(o"p�T�|�����G��m���i��$S`l�^|�E2�=0`�jx3w�Ӻ��.���� _�}���O� PJQ�;0ο��ߢ�?���/\��o�P"1�?w�Xr+
nIэ�C��YpO�g I7U�CxLzL#`ހ��Dk�K��x�[wL��h~���;<�͌x����~�j�G}��<DSW���Z�K���ׯ_?�]|W��H�6��IJ�Șb�7�x�/�S���xb�������:R-V�5��U��|��	���mo�t
�^�-� ٰa��N��K��hW���BOS��!�C۷o?B �9d�Ν;9s���Uu���=d�n�&�������x	J"�M��;�K��mLCu&�� 	TS,,�z5�@���ǤeY��~�l��*��Q�N��!y�ózF�/�w�M�qUA����#�Wop=�Q�\%��_�\_.��x%%q� �N��4���0�P���;���3A����(;Be�^[C0�m�_�?��m�ߠ���/(q� �P�����E��k�?!K���wI�ek��;��Ư��P���xA��(?G���h�)�#D�M^;�;aK@8��Sn��^��h�b��ⶐ�}~]�eyh� 0h�~)�����fV�����r�N�1<�.�\�R�r6w�i(O܋}'�(l� fP��ghh k/����#D�9���a/2���0�i��Ly���ۤ��i�?AYcp?��-y���g,�DH0�)�F�\ AC���_6�����BuVch�<w�K}_ $�r��l�G�L��d�1�b�����u�Z�b��?l}j%=�?2��Ca�7��B5�D��3�<#�x�	������-۾Q������Ai�h@1���h$���(/�z㴀�{LUԵ)����o��C�O&n��;T׏���=!q�*PN�)(�����h�����G�F��+&��������"�)u����6�A(�(l�}�0#��nQHJD@`� �%����^�e�\�hP�dP�~�ԱGyD��M^�5�z9�Y���t�ե=)5l+��"�nR�v%, 0Jeū�9qt�.��Q|��p�`^�dA�"z�5n���m��d�c�=���S�t�ɋ/�������JH@`p%;e��)bҐL�V\D�&�>���{"zzW^�KJ�m��O���~�m��m ��CJ�5��qLp�ѹ��Ы�9�+�N��������3�֧3�v��%l�����Yؠ�j��uy��e�8@40�8�]�����
��-�@8�i��f��/E��k� Y#�r,��u�B���S�J^�"lUr��@��(�
s�'l�oV}oξ幜C��k;m�-���ʗm9�"(xTC������p�?
���P��8�7ܐn28�j0lt���%�C�Y���g��5 t��8�}�����C%]Ј��aN
�&���D�0�O����I5L)q�j�&׭�< �<�A�c�a~�Eqq��5u٨��:©�
��l�A�'�s*�ݦ&A\PhS6�)hI��=�4��\�C:(B�����%]mp��L�H\�'w�`��r�۴ô~(T����A�2��m!Ϲ(ĪG��o{%�	�ø�ް�2�;�{<��C�a�8Ki�s���
�쯢�/�Vސ�	���Q@o|���̴���]���@̰����wĺnw9�m����T� �s�\˕w9����{�+@����$SѣL�c��3�&����ã�ئ�B�~Sr��W��,܉�g��$]^hB?�!m@��쳣��"a��h��z/E��^�Ʒ,�鹲mGb��s�B�F�;�r��G�za��3��7����i����^.D�u���Ƕ��M����C	���z�D�ɓ�t�E���U,08�db��:ݖUxx?&69��s�����ɢhfo_S?�QZ���9&�'�:M��RB��̹��% ��Cu#��d3�3�{2�ӓ�"5P8
�C7@�'�?�S��)��{�H��s&�N2i[�d�t�@�%1wo�mx����ݲ�R�P���|�I5ZM���lw5MJ��=���~�U'��v_"#2�c�_p�\� )F�H"�~3�$���u���v    IEND�B`�PK   �c7YuS3��  �  /   images/df606f07-93da-4db2-841e-5903537c99b1.png��PNG

   IHDR   d   2   �5~�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  uIDATx��	�TՕƿ�z�7�}h�D�L4j4b�ь:FL�ј��8�1F3f�q�*IF�b�h4��#(k��F/�[U�����(
�3��ޯ�߻�z�;�w�=�p�ؾ7H�D��x\�hW"�A)=]��T��`�O��JѨ�����l8�<��a�c$G"!��QX����
��>�={+�_`�d(*�$��^���xo�ڗ,Tl�2%���H�����@ � CV�q')|�$u�)�ޡ�;T_W����jmiQ̬1�ed(7/Oy��(w��N�(\_�؂7�2g�:�zMj�*���W����0�y����\%F����I�֭�ڗ^�{ｧu�}��Rg�466��z�衬�,�2���4���G�����S����_Wh�J5��~�?7[��6C0m�~�N�$���~��@8b�1����hmQp�(�\x�&�b�6-{�9͟���y�m޼YMMM***r�.((�֭[���l!#��o۶M555���������}�j	5n�z^u�2O>C�����１�A�O�a ��6���W��,�v��V��:	̗y��A���<W��]��h���9=��3�|m߾�� ����9k`�����Vuu���H�@���_]�ص �c�ѸCQ�{~�և�Q���+�ё��a�-v����/Q����������
)�Ԡ��g+Vc�D����0Ɩ��K��l�r=��l=��3ڸq�9���<����c���j3�����={����Y��6�g.n��w�}W�}��>������X���d�����Vǲ�:O9���>M^W[N�Z�2�)�|j���^}�����j�?��	
46�@y�ݥ���Z���4s�L����!L��ݻ���@����Z�h��*F����� �F�,Y�u+�f��H��Y�F��v��2E�w�T�E�W`[�ǂ.~�����#Tg�]��L�����-#�ѻ��:�`�t�Eʽ����jl���)���\���5X�xe�\�{����\@&V ���V#pQh9  \�V��W�Y�Y����P�M�,�b ������XNN����o��b�9�W�Z�n�����Օ��ΊΘ|��5瞪��o�c'k��^
A��z��Y���Ejʊ5���ʅ*��1e��4��RR:4(�{��;��g6��$��9Wݨ���7g���.�ȑ#��qG��Y�l�`�z�r�!h��ʕ+] �2�߭[72Ĺ3 شi��>�����V�f�r�8f�T�_{�v����ZwRl\V$n�����:0����X|���g{��@(qC,:f�A�*\�Y+�&� ��Ȑ=٩!U�$�4�G�H�D?_p&��.U����Θ�lx7�5��2����O��:���S\�W�?^�_��k.K�*�#� ��+��T_�_��{"�Lkm;�5���� �{]�b�����o��@�x��K�/��B3Ö�<���g��;����%
�߆�E�zB�vL��#t��J������?��	�<����~�6������\A}�������jM�qO�Y�������ի���wY|�߿���k����K8��V����SOU��j��',�Lb  jʹ��	�f)�h�jˀ^۳�V8�	��"L��NUd����Q���6f�ڗ-vV9���P��j3�̾������+5������Q��?Ӧm�����.@C]sss�;���^R6` X�� QQQ����$ 3��`�s���� ��z����f�p���Tg�����A�E)=ڪ(o@�������
�TPU[Қ�>�b�2�[b���ÏR��I��c5�}�V�a�%H�L(�3�p��EJ�|����Y�Ǡ��nT������Fm�UII��[�lqs�������wV�Ex�K|�Iq�c��"h\�# �]��Y݆\����5�%(5�c�/������Uv��<�����
�2�yH�n�s]����%�Rh��"H��-#�x8�=��A۪��08������S�2||�N1�o��+~p��Re +M��g�v�	�bx�B>�CHX���a#`c��<����+..v.+( a..��X��.^�XO=��;V��jy��ҖMƣ
�ۃC�E����*�����;+��gn�F�_V,���:��닕n�6���bU[�p����7�>�k�Bpc��<��R�s]���e�z��E%jy��O-|�Y���+ZT���>��4A����  ����`EX���_��o@@�A6X�O+�Z�8p����ְ���1\�8Y�;�W��o���M�����Ͼ��˵iPobJ>��xk��!�T��R��q���}�r���iz�nu�]���nR������<f��������n�g��v�I��u�1�=+���h$\�<��oi�	~޼yN�X��@'�m��aCG�\�ʰ K0F���<����	4� �����q������K��c(sqi��k�׈�L�fާp�9ߪ���y*���s4|����=�df�|$��ٱ/2��~��zڷ��u4�оt��N�Z2~�V` �0�����B"1�G������~Gp�H��{/�脊�;*��u|�]ah0��D�2Z�9lh?�^�>�3�}~�?�ߗ! P��2����Щ'*<n�����P��t����ߪ��#��T^k�[q3�����-nT}s��Q�,0z��Ը��@��m�� ����0+�X��'�&#!+�-w�ۗ��|���)n̗> �9���q�!r�Db�K�;�q_Çw�dO��q����H"
 �r!?��ڽ�}��8Ja|�{OeX��'��.'\i����;�:�e�Y5=��Gk0�Z����0ˌ�9P��լ߰�B�@p���ډV3�K!o oE^�9�ީT �����}aU��|�.֩����z_��T[�R<� S���:
~q�:֭UÕ?V4?G#�A���UT��xr�O�U����M��Hf�_�ӳ84R�}K�����p�СC�`����!,M��X�14����]b��<��瘧�)���20���+Žm���w�a
�=9���Y����_������ac՜�嬃�v�`�z��ʟM�~�
n}@qKb�'RS�/Ġ�`l.�_��%+\�F >Qcc L�@ (���p?�m!p�aŊn����>>}&���s�ǰ� v�Ԯk-�,~cEI�J�xÎ�&�[u%�Z8e��MK"��K,�m��e���8�oZĨ��/��H�؉���'As��"^G,+���#ׯ@�#��a��a��(�WW�Fs)g x �
p%h( ���ǚpUX��s��W}B�'�����qM� q��V�B�1�[��9܋����a�`A}0b��L�����r��5��$p�6sy*<��H�&�8L�Go�[���W^��3
���y�;�1��&�ܤV�6oH�V �*���Zd���\�� h:��ԯ_?WF'� _wJeb ��0�r��B����<ϼ8��qy��J����u@P�`�a���u%�X$������'nk�ˎ�=��EkG~��ڍ?1���(�-ا���G�:�3t�ʥ���骽�\���#q�$я��~���n�w�H"��I�@��ݝ6���F�!(4��G��Zܕ�<�e�{6;��6�q�����P�S��~l�1?��o�>�z�	]'I-N$v��D�%G&)�e��N9�e�
c����T������;֮R��iʛ~�r��#5��1�k�w����j&\�7�â�Ԓ|ل	���(@�WE� <>�"8J��qV��C��6s}b��%�B�e�c�Ǡ��ꔇ$�S~u�j��Rr�n.k..�9'K�֬;5�3ץ��z���h{�5WB)��_���e�N��R�L���	�jy���0�,,R�������� >��~=A�}������O����b)9Ԯs������3��z�^����ۉB����׀ekT1�/A�����7,;�c�W,�v�1����Wn�%K�k�i��[�W�k/)�h��!V�U�'S���D#Z�p�8b�s��G����o`_-�Z,$q��䚶���U@�������Đ�Z�/s%��ĐX�j�*G��O�֕��N���Xl�����$xwu�W���.b�zn���.-����[���2���~T�54bޛJ�8�����<�d\u�+���۶E�>�������IS$ۏ��y�	���k���w1Ā�WW)h(줯�@��à���|b�C��x���#h0�8�[|c����Sg>90�l����z_��$8�]Rls�TU�x�\��40���"��P1��K#����]��&����ល�4�^5?1Si���@f���8+��ť��+���J2����Ծt��V1�%jk\�@�K���BKM����!3?51D��a���A�������Pq9~�
��C��=|�į�@ �R�-�X47�X�2\s�4�z�rq�����,^�EM�����_ݡ��np��@N���x��qB�Wy��dqѬ%:翓׈w��y��6)��J��=�U��ofcc L���g�Ԁ!������V�db$>�(�9 ��X��]�$���!�c9�Tf�1���Yيo�Pˋ�*��8��V��@��ؑP��G��U���?캣v��Y;�7,�S�a�#ʱ��G7".�����y�O�c9�&��!�Nn�'p$�>1d`��>1�ڞs�9>1�X 3b������g,S�����}��T��3�-���I)�K�w߬Pi7��Q՜��Q.	�5�����[% ����!�|��X�K�vZ����I������KMqO܇�y��o�%r|�������s)�r��l�;x�6ZVޖ���A����,�)�`��+��-6��{.	W�c��� �V���8�3����ZXڏE� ���pE�H���C�X�3Gc�k�YH���X�ɍr�P0��WY���h�F�l��L6!�5�&�x����4��}<`��Y����ɚ4�P�P��xx�ӯ��	�w��@h�0(�we�c�����`m�N�G��\B߄P���ۛ<y����̼[�<��h�[₺˴;��@Ff2�|@c��~��5��`A>�S�x]m���-�� �LV�,?�^�L��(�\W:����V#��D�@��.�b���XF:�5�~��t�s�=��p��µ؈q�:H[7���ٮz�׍r%v��i8A�]1��f�t��O?��ƻ���Bݕ��W��T�w?�-|S�W�D1#{J<�~_ ;'�dLx�/�Ř�5Y���{t�	'h钥�~�n`=��P(��������rJ%�9�9�_�e>�s��Ua1X!�+��UE�!���?�x�8@��^!�,���w4�u��3����;��,��{�q�E�-�(9F�n}й4����ܢ��?U�.S��:#�v���\m��8��xW;��J�M�\�أa��aA2���*?�`�t�T�u��N��R���ʳ-6OM���> �#�$���{|U7�Q�����5'N��	�����槞�Z���F9{ ��i��d�x�2�<Fm��Vd�r]XK�9�^�(�̟݋�4G�I�N)�h�q�����2?��ٚ���]�m��=4KGw�6%��(���s�zj��,L��a����@�2��^,�o����}A4N8�Du�6%��j�ۺ����Q.a��n�e�wJ��m��b�� ���]S����9Na<�YW��4�ۘ@OU�w��������r�ׁ@��x�G���Ć�x��4��SN=ձ Zv a�龼>�`x-���VR�5|)ē�~�:�QX
������u�)�h��#�|ݕ�/[�bp�OޫF9���Qj[����
�W�0x�Urs��C�HE3D�҅�X�J��~�k��8u.�w��KU�W?���2���R�Q���g��н��b����v��i���Q�z��m�`�ܔ��+v�m�?�9�|,!��_�@�~V��~����;f���{����,��#�	�4ʽ��:_��g���z�{a�ds��!�c�su���0\St��֟�_^�\Rڨ1�Ν��*��.n�Q�#�qu�OzG�kF����4ծ�V��ǟS�ߞӎ�ڙj(��-�ߡ��|���_�r`ۿ}E���H}?��m����P�<�����	�X�gV��=m����|�H\;��ϐl�;�<�zF�Q���5h�L��6K
I k�;]1J覥�d���Q~�^i��B���sg�T^k~t�+�8��O~R2�������'9*K�2���:�am{\#�XL����ʴ�1��+۴w��Oꭷ�vV��z���w:� �Isv�N҈k�:u��y��q@���KM��<�D�1��.+D��:C�����O�~amJ��52t� _������@����m���5+?�;��S��G0������B���~�Ҷl����|�؁���Z��'7H}?�����!X�?�K��͗K��L�<E�9E�����HO�Cw'崛����!3?�]��~�kѩ5��s{���df&���;j}��J?�+����K0R~oq�=>S��������o~SC-?xu�<���+N'� \PjP'���C|�*y@�ʨ9e�&~������`�"�2E�k�3�H=�߶x�'����u~�=T�5��<&2|Ծ�I���t���me�y�9�w�9�t�Z�`�cC��3:�j�U!l�	�a��C�E��z��q�?t��-�m����{�h���ԧ����/D��k-����;I����F�E�?�Ai��I���ua��ȯ��!����Tרb�m�l�]���-|)�D�X�%���ܢ��M����۟S�c�(�nM҅�ao���:A1\bh�V��pQ�S�m9p>���Z[��b˵���~�
�͒�� ��V+��h�Z:�W�߂�	�t.�f��0��S|������_���[�^e�"u|!q��s�L\{��*���Ͼ��/���f��'���7@�C�g�UAiY����f���Xd�b׫e�j�ֽ��M��Q��/. �2������+wfw�倒[�uW6p���o}Xp�������Q�1�C�I��� RIr �nsI    IEND�B`�PK   �j7Y͆F<,  �%     jsons/user_defined.json��n�:�o!����oP��:k��vՑ�jr��	ɪi���9�t�%8u��/��8y��5�=�M����˥�?G&NR��o&_&Yj��=�,���e�����\ͫ{ߟLG��Y��>$��ҩY�<Y�����D�c	#0��
T��
��S�<2
靽/����a.�4�!�D2cT��V�����6��EY,ʢ;XU7]7��li�E���q���>�u�i�	���U�'6��*�B�Ňl�TŜ%3{�!���~�W�4r\�DC.�U9�q�ﳼ�Q��6��
MuCn����>�L��`>ȑ�WB��g�����,�-'�?'���]nL�bG��I��H���Yi�9�A���i�\����l��D�do�t�=TMt�0Z5ٱx]#9Ͼ�pV��_����E��o�첮����}ߔM��9y\��p8� R�&�K�����"=���:*Fn�eR�ܜ���2�+h�qZu�+�J�X��M�4���$O������>Mt����C��!@�S@�@@B�@��CAp ��?�^d�I����!�4Ww�}f��ڟf���V��Q�-��,�e��;3QK���ڢ�N��R@j`L1`�):�L�ڣ�DYS�&GC�
9a@K��q`�^��� ��c�Z(����l.���y��r&;��T�~L����ee���G=~T�͖l��0���;T����՝It��;{�'8U��O��l2Q��n_g3�?��go�A�yU�v�ǫSv���VG�ϸz��j��!�i�l��yh��Eܛ�4ZnsbO�6�^��9B@�422 f!����"�!(0�App��#�����yT&i�;���;���������ȕ_ Nt���P"BH �"��}B����T2!@0��� cd���C����kX)�������Һ�'�ѠB<R�dC����v�Y<��Z�1�1�):����A\�+��/L�ѥ;n�@=#\�\�\��c\�g�w�S�>m�Ǿ}���E���<o�����)/���W�9��z�Ν�ҭ.|Յ�x����n�t�ɕn�n}���.p�P�������Sw�t��E�������	0�p�07���M�yw�n�8�Ę��M�&̼�Q�w�&ϼ�S��D�&Ѽ�W�݆��L��n=v�)nR�;���=�&ռ�c�ݓn�;{��=�6�}Q�l��d_��nW�m�b<�<y��F�/���+n��ߴ�����G�&�t�@��L���0�3L��&��W�x���T��e�8[�&ܸ{1/����M���8y2~��W�,۽�������Ve��n����ٮec
r@Zm�1B"�a(�8@氏y��<�c�1�>��B�_ޖi�dft���w�h[���Mr��de�c�{�2u����Eh�9�& HhL$���J�PĊ�����H� ���`�����*��E�.i���·{~��4u��$Ci��]�xY���q��ˍ:v�w���l�l䉧����5����@)9�?&����=�9�1@�HU���J�LB�R������/PK
   �j7Y#
���$  �c                  cirkitFile.jsonPK
   �c7Y�/WYp � /             �$  images/0f73fddc-80bd-46e2-8805-d6b40fad9a5d.pngPK
   �a7YmS�;F� � /             �� images/45855a06-4846-4a51-b2b1-60b9838f281e.pngPK
   �a7YN�v4	� m� /             2> images/4949577a-1080-4c93-a0f7-9bc81c12f32a.pngPK
   �c7Yd��  �   /             ��	 images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �c7Y�]��N � /             �
 images/907530ff-a8af-4c9a-ad67-f4101e76dea0.pngPK
   �c7Y	��#u } /             �e images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �c7Y�h�F  A  /             G� images/cb0ca54b-1964-4771-904a-f612fb73280a.pngPK
   �c7YuS3��  �  /             �� images/df606f07-93da-4db2-841e-5903537c99b1.pngPK
   �j7Y͆F<,  �%                jsons/user_defined.jsonPK    
 
 j  u   