PK   %:Y��+%  �g    cirkitFile.json��n�ؑ�_�� �.�TN�/�o<�������?l�`�2�ܭ�ZsY��/�ϴ��K�dK��x�� �c�������<���]�}�)��-�ow7��fqIa�x[���?5���zS��w������=�;��t�&�][5�mS���L��o�*�+�&U��ě4䔇��Ҕfq�����
$V0%��
��b��)��A�`J/f�*�2��
�L�RSfb��)s1�T����A�k��P�%"�T�k%ɋ�X"R�˥X"R��X"R�K�X"Rȋf/q/p����%�j}5]���^U����8�f!�#y	�%D{���Ѧ�N�G�.����K���0�V~JKD
�)A,) �g�)��O	b�H!?%�%"��� ���S�X"R�˸X"R�K�X"R�K�X"Z]y�KD
y�KD
y�KD
':�F�N��)�;�;a�;!��.g6Q@����.�¥�4�f��T~s�s�X"R��ab�H!?��%L���0�D������B~KD
��_,) ���g/���%"�|�/����)�����KHN�>G^��:,��ggy�%$qy�.�p��� ?%+�	/�	�%H]Q��	wB~B
��X"R n��OHA~BKD
�	I,a�
��"}?��������L�� �D��{�D��{����3�)��D(��w�a�Kg� 4v�����t����Yl�t����%l�6vP:��E/�����JGX�8���.`c�#,]<�cc�bc�#,�)3l�2l�t��3e��]�����t�,��+������O����G`>~�?��@��� �� ��������2�|�����;,���Q}p��n�G`>3x���߀Oty����~�g9]� ?ص�D�3N^�?��`���O��{,��x���6��`��ǫu���,��x�8~��+�,`�c��ǂ����|��?������W���v?X>��z:p����G`>^	�ؾ`���k���,��x�%8~`���#0�?"�X>��Wp����G`>^���`�����C?�~��?�8������&#� ��I.7�����@��/l_�|��E��������|�|?�}����ރ��/X>�q� l�<ؾ`�������,���M8~`���#07� �l_�|���������ש����/X>�q;p����G`>n���`��g�W�z���$�|.����=�W?ؾ`��g���@J���o��G�p��`����G`>�H���`���͐���,���8~`���#0w���P�R�~���������v��v?X>�q�1p����G`>nu�ؾ`���Mڰ�K���G`>n/��`��Ǎ����,=�Wo�]o7�f_6��+�B�%>-�\��$k�k�.���׌�~��p���~�3���p�9������]Sg?mw:s�i�ҙ�O{��~��sn�H�N�w��$�/̼��	������s��o𮻹��7xA���Һ'̿�������fs��o�ڰ���7xU���0��ǚ;^z����uNs��o����o�������J|���$,�I�l�,k}n�5M~��M~��M~���ժ�����2'�q�Y��%�OS�֦K��}�4��}w��p�$qk�Ҥ(�"��ug�"�X�?��&�ϻ:)��b޸<���;!�Җ����y��'?�顨C�l���8��ڪK�,O��|]���}�p᧟ϺI��gݤ�}��Џ/�۲�^mw���Ͽq؇s���'y����#�!	�C��C�SC2�L1D !�fC2�1D !ÖC2��1D !�_8 �H\�ƕmX�&X�F)���	�	V�	V�QJ���b��o����_ �`%��Dy��K/d�q���/���z�"�*�V�QJ���b�ͿqpX��:�R2�M��[XG)���+�	6��:�R2�b��[XG)��B6Ȏ�긃�q���/���pWR�o�\!d��qw����+2���+�����F��k��B&Xw�:�R�N0&Xw�:�R�����:�au��+�aL�:�a�q�� �1�긇��QJ�����V�QJ�"Ɣ���V�QJ��v�Ǡ��B�3����gX5��:`u����`L�:`u���`L�:`u����`u��k``7�a��6G)�Z����GN��U�EURa%VS�.C����J*��<]�W�U��TXMy�6�
��+��Fߥ�Ӧ
�h��
k������&����(*q=m��+����-\WVRa5�i��*0����j��6pU`\5XI���	�1:�K��th��f��*�.%ۥ�H�x���R�%Z~�\'�:�K��th��y���80Zҡ�g�ub���ThI���0��Vǉ��oZ�d���1c���Thi�vx��A�1d���ThI������VǕ�В-��ѹ����ThI���*��VǗ�В-��҉��1�[b:����2���ThI������VǗ�В-��Ӊ��/S�%Z^��[_�BK:���R'�:�L��thy��Nlu|�
-���ZW����2Zҡ�5�:&��2Zҡ��:���e*��C�k�ub���ThI��ׂ��V�iE��u|���eNǗ�В-��׉��/�E��Q��:���e*��C˽tb���ThI��{>��VǗ�В-��Љ��/S�%Z���[���ThI��{���VǗ�В-�Dщ��/S�%Z��[_�BK:�ܣF'�J+ɔ����2��˼�/S�%Z��[_�BK:���H'�:�L��th���Nlu|�-�Z�
-��҉��/S�%Z۠��Thi��ls��eAǗ�В-�8Ӊ��/S�%Z�զ[_�BK:��sN'�:�L��th�w�Nl��|(����eAǗ_�BK:���P'�:�L��th�'�Nlu|�
-��roI����2Zҡ��*�Mu|�
-��r�O����2Zҡ垥:���e*�4�v�[��t���r�7�L�3�d羧�r���L�3��g���n=S�L?�*gzQ�T9��ynց����^�:W���^�:W���^�:W���^:W���^�9WT�1Y|�-�se0Y|�]�se0Y|se0Y|sϺ�,>����2��&�ϽVo�&�Ͻ��^��m��~�P�W���U���>��MC�e�����I*O�I*O�I*Ol�ZuTהUf�4=��+�$�ij��ti�=�I*O��ի�y��A��Ҥ(�"��ug�"3�MQy����yW'5YL;�'y�/	Q��T�&���,�T�d	EZg��X�G�X�U��Y�z�����2I��d�NRy2w'�<�Sz�r�-o�վ]\�����������磌�|�_9:=H�	"��!� D �C�B�@B���"���/@�@B��� !	��2�$d�K""��9\^��H\�ƕmX�&X�F)��U$�v�x������	V�	V�QJ�p����+�(%s�&�a��q��(%s�Z�a�ͿqpX��:�R2���&X��:�R2���&X��:�R2��&X��:�R2�K�;��V�QJ�p�Ä�������V�QJ�p����V�QJܴ���V�QJ�$���V�QJܔ���V�QJ�Ƅ�&��(��V�QJ�X���V�QJ�8���V�QJ�v�V�����x�+�	V�����x�%�	www{V�����xQ�	V�����x�	V�SXG)�����:~Ni���1��a�@�TXI�Ք��ahU`\5XI�Ք��ahU`\5XI�Ք�fhU`\5XI�5�.���t@"��J*�q��A�H4XI�5�QT�:����+���rМ�
��+���rИ�
��+���rД�
��+���3�:�@�q�В-?۬[%ץd�t|�/�q^*��C�Ϛ��V�}�В-?3�[�BK:���Nlu\�
-������81Zҡ�:��qc*��C�kJtb���ThI������VǕ�В-��ѹ����ThI���*��VǗ�В-��҉��1�[b:����2���ThI������VǗ�В-��Ӊ��/S�%Z^��[_�BK:���R'�:�L��thy��Nlu|�
-���ZW����2Zҡ�5�:&��2Zҡ��:���e*��C�k�ub���ThI��ׂ��V�iE��u|���eNǗ�В-��׉��/S�%Z�1�[_�BK:��+A'�:�L��th��Nlu|�
-��r�
����2Zҡ�*��:�L��th���Nlu|�
-��rO����2Zҡ��.:���e*��C�=jtb���Li)��/�:����2Zҡ�A:���e*��C˽�tb���ThI��{8��VǗ�В-��҉��/S�%Z۠��ThI��{���VǗ�В-�8Ӊ��/S�%Z�զ[_�BK:��sN'�:�L��th�w�Nl��|(����eAǗ_�BK:���P'�:�L��th�'�Nlu|�
-��roI����2Zҡ��*�Mu|�
-��r�O����2Zҡ垥:���e*�4�v�[��t���r�7�L�3�dg����=S�L��*gze�T9��z�ʙ~�3U�t���r���ܬ%/&{Ͻ�u�&ϽZu�&�Ͻ�t�&�Ͻ&t�&�Ͻ�s��c���[*��`��ܻ ��`�����`���{�u1Y|��se@S	L�{��\L�{yݽL��*��*�&���8M}R9��*�Z�ۧ'��T�<ܓT�<ړT�<�v�ꨮ))���iz��W>tI��Դ���4{:.�T����W��&��XťIQ�ER;��VEf�1���$��C��N
j��v.O��_�*m�jM�ɧY&�<��:��扱>�*��j�.��<�&�ua'�e�
���ܝ��d�NRyX�>,���q_�۫�\7?..������)����m�����v��|���3�F����po�"�c����}A�ψ"��U�R+ı��D�sڛO�#�f�vɓ�N� ��ߺ��O��>9�x1���1���b<���ғ�����	�QkN���pbR��y�k�m����jӌͣ^E�����?�߿$� a�{�:|��w*������_���o��a_9P���~y��H��X.I`��W& �?�!����j������\ё�^EF����
p����Nܡ\��e�CM���>�cB\=��M�����p�.F�Es��l˛}�o�����'��my�n��%I�w�K�X�p']H!�8܉R�%w�b�Ó B
����R�%L����B,a�Ƿ�b	�?�-�K���q!�X�?��-D�D�O@�$@�k���R@%@�k��3�R@%@!�5���y:*k�q��X�R+�0�UR�b��(�rsXv!�@L^�W@��+�0��#R@��+�0��+R�4���\�V�H9 ��ʫ\���H}'��:@=�k��
")�r��:3!���K�N�DW�� )�
C,#�BK�������t��P���'9�4;@i�k�� � ��J�\���8 ����rn�� _���5�)7�PO=���5��3�#���7j=���5��0�.��G��A ��/ �o���_ ��02MN��4@i�kp�Q �4@i�kpK �4@i#�Yxq5 J�\��
n�f�)`�+��vu �����y���8�C_;����g�A�E�$~X>�r�^�����|�����A��#0_�.������G`�8� �oЛ^��X>��y 8~��������ϔ�V�8=H��|�3堝<N?,����:(�$~X>���	4ځ�		M�O��cw!p��!�6"�v"`BB�Ӻ�����Є��1:�hG&$4!?%��!ڕ�		MhK᠂�O��W����Q�LH�fL8������ψ ھڿ�		Mȫ�1D{0!�	y	�26�ŀ		M��/�1D�0!�	y�:���)�*hc�.Ƣ]��Є�dC������c�v1`BB�R)t�.LHhB^慎!ڶ�		M�K��1D�0!�	yy:�h�&$4!/D?.��)`BB�Ft�>LHhBsԔC�O���w����/��_h���>š}
��Єf�q*�����*���>�W�C��-`BB�htѶLHhB^���!ڶ�		M�K��1D�0!�	y�<8�m[���&�%���m��Єܮ C�m��[-�c��-`BBr�t��V��Vжţm�G�0!�	�=:�h�&$4!�A��S���&4���A11>ցE��	)ڶx�m���u�8m[���M>�J�@���v1`BBr�t�.LHhBnR��!�ŀ		M���1D�0!�	�:�����h�.&�]��Є܅C����;��c�v1`BBr�3tѶLHhBn��a��-`BBr�9t�>LHhBn���!ڧ�	�)�z��z�i7��)l^Q���(�i��%Yc\[t��6��q��A�Ù��	g�tm�9~�mu��A�ԙ��Mg�t%�9~Бt��A�Ϲ�#N@i�A7W@��÷���f��]ms�y8|w�\i&_6W@\��8|��\i&�]5W@��÷E��f���Ls�i�L�i����,�����
H3q���{�ʷUZ�UBM^%>�Wq����r6U��>��M�&�� N��1�4��ChW��Ꚓ��L���Yj�C�d>MM[�.M��������ի�y���y�K�����v.ԝ��F^v>s�#�o��������,&�˓<���*m�jMܥ�>��G>?uh��c}B�c�V]Rgy�M���>����K?����4����4�PA>,���M�ߖQ0����)e`q�j����w�/�o���4�8�_�������o�o�[oJ�-���[oN�=� ��G�^�GXay���GXay���G8�z�x���f�Y.�|���N�Z��O��=:0%�L9����M<��i�|�˸!3�>U�̱g�+��ǐ�
	�p����!�R&#<�!5$4BB'�v��h�|�����=LE{ؿ�G�G��J�V��݋C�L
%|�s#P��K.z	L���!T8�z��2�e}�2�5}���/��U{ť}X�j�/�@�i�+;�������������*��������*�*��U>�U��U�iMuuU>��z�m˫�͞�٤�����w�m���x�_�x{q�/�n���='�'�Џ����W�*~���G_���n�n�ݻ���	#u�߭7��(n�w�o��r�}uu���ϗ���o/S�{�ؼ�q�Y�Y��w�v��W���,.��ꦍ��iwY߬WW�ǟ�ڿݮwm�����c���vU��ݵ��Hn� ��/^�;��@q�wn�_ocP^e���-mf/��-ϳ�oF�2�~�u'|�$���wq>����n��,�B�V���xT���n���"N��զ>M��.��:�T���5k�w�U{w�_�Yv��]0o������k��vl�7���u��v۬��fA���o�X�}�ެ{��P7�[>&������'�w�������;=���u�M��.
�2�"�*
|�MQ��?o���)ODn�?l�
��cp����������_����o���?�o��9����şn߭�݋��/�Ms�(��(� �2,�I��M��w&�d���K�63�5�ZW�"{�U�l���dUU.1�͒����:�:�C5�0�-�~���0��i��"����L���SZd�[�y~��)�$�$g?1������ß?7��L>��z}���g��v������zX��O���RW7U^'m[��wY��+��YcV��Oͤ��tnZ��|����')��7����ij�X͎o�F�{��X�n5�Ml�S��������IZ~��;����IZf
�0y|~��O��͆�3��0yF7$��V���j�<�[�gl�a�n5H�ѭ�3�� yF�$��V���j�<c[�^��a,��h+�j�5,�cZc[��$����+�Db���Io��Lp�n{մ�����9��������~�z�|�X7�O:W�S��$���x"�C͢M���:di�A�۷?^_m�����﮾<��4N��%Mh��$*�8�^%MSPhW6�K�����嶳�]5InҚ'*.���USQ���8��8�������`�ũLn(�Sg9u�&+-����dyUԝ;��͗�oZ��c������{����U�PٸU����y�D"׸���M���P|^�v��W���J�f��.q���.lRx��t��:�+ߌ�|~��iҬ��vf�&L�ڤ����kr�eիp����:Nd�8���a��}�զW���e���rSm���[���4y������gM�kon�~�a�g�[_�#�u�����0S�Y�;ɉ�T�jc@�z-XS�غ-�fX�99�&���1����є��(rc�2lUuE�u6IW&�8�N�B�bG?c�4�;�a�jL�ŉP�}��lU$E�$�������<<���?_/�߮�7����_����ׯ7/^��w/�ǽ�i{�;��o��m�k�/����͋m��]ƭ��>�ꅮ��q�w�z3"�k��j�6W?=;��^���ϙ����,���|I��G�.���WO���ic��p��EK��4��8k�8=��)W���n�Os'#W/{K;�󿇥��8��٦�v����/7�-�io�޶��Ej�c��_���/}�=+k�U^�IմyB��It�|ѺH��X��I�3�Ʌ	���!����)N&���l��lOc�?��|h{�sa�^�����9Ǐ�\�C�v���f�6��Hӏ?{��ߖ˅��i��=�O�t����T�۶y��.�׻v���/�����i�W��|����<��/�`����n��zsw�=�q�7l�9�c ������'y���U>����P��ޮ7�����^<N^/�F�W����o�
q�?�|���2�C�,ǶJ��Vo>�)bL������'@0�8y�F/��`~n���d��t��cPM����� ~�C'���8>�Ŕ:�n/Ƕ�� *� �	p�^��W�1��	p|+�\8�j�)@!��	��|R8�f�1�pO���ӭ´o�i}]��{��g.��:�}7'��~|��?������L�=g�|Z��6�]�&O�M��<�b��%�񵒳�"��Gw¦n51y�	�+����C������Yy�SM6--�s���<E�*�S)��+���)s"p����\g�8����#[��	=v�?ǯx�Sk:?7�'�rl�3΄/�������X��ݺ��01'n����m�Xmn����w_��w|���Λ�����z����ޭ��/>�?PK   �a7YmS�;F� � /   images/45855a06-4846-4a51-b2b1-60b9838f281e.png��eP\m�&�2�'@���'������!��Np������w������TMͩ9��i���EyItTbTti)�2<9�2"��[$�����3̡����O�#������������)������'c{ۼ�:�0���b����v.0b�vn�N.�&��.��{,���$��=9�r��5Ɖ�~���U,��u������Y�|���ڳ�-��]{&�I��<XT���2_XT����!�H�k��H��)�E"�]{��P�$K�t�u��t�A�(�+=�x�j����� xK
�2~�&�w9�b�]JY,��nV��7E n4�<�:�1�я�������#������ؗ�3�\)�0SJ�6}�5 �!0���E��Vz��|�f��@��'��c�p:߷��T-�m�������ru��� �d���1j�+�>ŭ�3��!�/{�h�1B�0�m��R��L~�_B,�Ik�li]�(�:D"J(k$�6(O���x��HL��MZ4�4A�B`!t}�>YZ�Ț? �Q�@�Dy�Q�ۭRV�P��>)�Lgq薰�MA���@:�7��B���x Փ��a�Ӂ��Y�o�zϱ�(C�Z�潀�gB�P@�L?�h���׸3�î���w��������2���kr%���>��Z%T��ǂ6F�G����Q�!�����+c�#+�VC�	[�8�>'�C'�w�!�P�q��5�6�7�#�(iTšq������BE���/ Ȇ����uvB��a
��{��b�����@~��X�R�p�p#>�\�mR����P�4�J�G�w����� �ԥ�]�X�D�/�-]h�͌C�TR����.	1 �X�qw���޸��~��tC��Q�S�&Fۂ�1\��b-w�9Y�����Y*�U�e���C�N�X4Uj�Iړl�{���䩋�{�qSĊ]qm��K�Q.�2���r� B<�6
;{�55��G�� ��M�8(����@�:��ݎ�k���-�ŭ{=`>�.a�vtVk��\�_:��ȷ3�w�'���#RQ��`mlx�3
h�8���t�$#��4���=I2t#�S�t��Z&�
bK�@�L��
|���F�8<R�(�R������j	:���٪��Y-oߏ{ƍ&�]��%��Rţ�n������c�:~柔���΋��g=)/�v��j�0�\��	{$7�:0�H�c��lx'���o�MVH<�m�ɽH��5���?��S��p�m��y[�o�]����aa"��A�^t�S�.������w�v�,'W�E�`l���7c7z�G;����r� j7�m���X9�Z�1� �Q96����ϼ�ة�ߓH��t�����>��ml�s��Љ����&���|ɿG"6D;��̧Zl��yZNY/{����I&�}vcD�N&AM���D@�5p*�e����*����t�oJwz�)g�g/��_�b<��7�$>M~舙�6�0��I�\��;Q(�*�Z�M4��6��i����?�%�/�Hl�X@�L3�ɸdSO���<N6C5v̈́�޽���w�!�����T�uJ�0����-Ń�-��*L�c<"v�����W꾡���� [��G�e���Ň0�~���sw(������#�l퓔��\��z=[@ؙ��K7;�Fλ�#�0��������:B�����b����ο&L�)�D�,�1�}�"�C�~(i��M�Ƞ��Ιf��#)��0|��K��KBJK�)R��`���Z���?+B�-�����fI���0�1Wa���H�N�D2��	i�b�嘳�fKބUvK1q�������{�� �]Tj�<l߃R��-�|R�ИLBQ�eK�"��8n�]/go8�,�L�Z*F���ec*��"lP��>f�3�1�N��Rz`߫3�/ܝ��Sq0�4�=�F5�!��ĢP�}���f���%��x�*����)�?v�x[�����6���J�����|b�>�ّM��K�r���O�2/�	&�ߡ���I�������(�r+O�3��;�_]byU�dF��A�1 �r�����i�-_�Wn�F6��N6����E��\��l!��9�޼{AP�_����z&y2�_Z	V��7��	;�w���a
�[N���p�k=�d�%4�A�1Q�k��2�%I)"���g�͍z�%��fc#�ç�
�p;��!qȷ�|�5�w�҉9�=H�@������<��R�Zˈ��	ʔӎ��0U�'?���%g^]��y���P�*le6�R���I.O�����B�~����AIY*��I�۞T9�q���u��h�+z犯/��hI���w�[1gu�S=/.��[r����M�$	�V��J��5�TC�����q�*]^���Lv]����6�˱�h'�l�`/P����|�!;����6�$+�v?IFZ�܍�/���j&��x���b)��O�D��v�YWiY�>�+�2�b���:����/��wA���v�q��
�Bg����U8���I���_��`��~����y�|���k�P�֎��X�y���.��ږ*����wp�)��.<�� I.�l�D3�C̫���4�H�3�|
C�����l>���@��Ћ���7�Ǵ78�D+����B�[�j��0�����2q�U��.��ƕ�&��v���|��u�ʁ�J�Ձ��(�J'28;��Ȼ�ђ�]Fq�>}vD,�J�z�G�ᮅ�I>C��0��JW�E6aߩ�yK�e���>*7��W�l/R�B�{�;�G�r������_FutG�y�����p�DR��Ä�8�0��-S"�m+�M�io��w���H�8G�����<�������T/���@Q���,
�[�T��>K�ܯ=��1��L���[!�P4JS�c�ʔ��-��ia��E.��ߋ+�ȆiW�|��n��;�܄H�<�؜O�N��q-��GAQ0C���u��y�F6n��3_�Eo"�&�T��|"G�.xC?s�G�Gs9r�z�-�߭�z*qg�\(&�l~�pd-��ߺ��H�����x|��SH�uz�S�䊠����Zj���5�aL������2��G�`X?�s
�̛�Ž+To|�����:"�qf�كkH2|�"���*��D�����ը-b���QQI��[��l�Ae��	���� �!(����M�CUj�A�4�f}���
L^�f��tݱ�B�������䀁ǌ��a�Ʒ�\��u8��{��4��_�]���/�6�-DX������r~}yw�v�y�/��btěhFZ#17ф�nPo��/�=���mX�j'�n ��%k��OZ3��0W��/�癴�M�X�b�tvK�8q?� ��1:���Ɯ�`6��q�p�صN$��R�y���e����C��2�����'��ҕJ]֕�S7R�Mxo�|���md0�~^h�9�}2�e6t�5���L�Sö��Z�a�NI�SF�S��o�bt��`,T��o<Wұs���a�������RL)��SQf��dGz���\^�sf������6p�h�4y2���1��5D�p�6�hl�a�@9���y<����=14�� ������֋�N
y7z'���C��R�#Qxb2Țˮ�ב2�0F
���?�� d�o8�.c�M��׵%�Cey��a�8uU��z캛�ω��MlR9��r.&`�%�R����4|h4�jN��nLCc�I>O�;Ϗ��,����i�,E�C��31g��C�`��=D�!���Yg�M���j+�!��F֔���Thv��90f{�Μ+���s=C�����}B��9��wyT�K&y���a����8��-�ӥ�U�v!$%����2�4��!�,���%��-����k���W;՘fb+$��<�d3�8�ѠK 6�� �l�f�m�Л����%0ɢ݋7Ѥ�V�y��D�x�~���f�A!;�����
 PD�%�x\֝��&GV��9z�R�\S�H\��94>lz'�ec��޳���2A	W�r���)4Ht����X�j�����6\H����nH���6#�,��6��-u@uLj���8�$���f��f�b��o�$���Z�<1�����a�Ҹ���A?U*"�ݸm���6f��M_>�eE'�%���;l�~/�2�%�0P�I���)��ۼ�6�Dm��;�|�,�CD�-+���<��w^��񖁴��Z�f��``���(�3K�ߙ+b6F�Q2vB���_��]��P�f��X�����m��9j7�����m�6ǀ��4�ǉ��{(|�hUK7���eCl�6�^?F�[^��@���c���#���C6��R�#�V�N!��fȗ%�qO��������� ?��P�����bn����	K�2T���Qt� U'�-6��ÇQ��r[�D�3�n�>���q�?�]����t&��Gs̏�B@����=�����g������+Ġ������$�m�-:������_L�q!S��cݶ촛��>hPR��S���з��l�z��說r�j�\�k�Du�p���s�[� ���J�g�2y�t ԭ��{L�cޅ/����gFb_����ʟ�sy��<���N��[FI�R��|?���4wn���(`pccx(3O����B�@@z��P�ئ��7�Ɔj��z݀[%��]�*��yg+����+N����>+��kx���H����
O���e>\:��B)!Z�ߧ�;�x{{ >u��������M[
Bg7~�w��0X��LF0е��5�>̣�SB��7Y�����pJ�Q��ʵ�]��p���V�,1کx�^Mk��bz����m�O���,Zu�09I]��j����Yz7�[��4S"+s��I��W��4�S�UMܲx��n�`�YԐh9����+����<͛�=�C�]vL@%��B֩�w$?�jq0��{�
0"���y�����8�JCJ����4�\V%��
�Ɨ~��\yfpB�l����^�gN[�8J��}w��Ī�C,a�n#"r��O���4����\��7�v꿉��ゎ�r%y���q���Z����x�漀�*�_.B�b.�����NG{,_ �cq���2���%\��6U:+,cm>b?����(I����Dp[
�wk���</�o��n��(�1GW���8PQ����gxIB���7�tut/�S���6?=���t>�i)�.&Zƒ�G�������j/��"�2t��^�����qG_���#�HؔAkZ�^	���DO�(I�~ҽ��m��)?/����b(�����2����ц��&��1��%�4I>ϛ.������P�^�Іȭ��G�s��Cm�lO���n6�(�v½���tO��#?!�V�$3�'�����Ψ��줨�W����4��S�֙�Ht(Qs1m�I.T�0��P�������r阒B3D�^1�s���ح�x'k�מ|�yRt؊�P�\����/������ti7�fbΗ���m����U��/�v�\ԓk�a�\>�|����L�D̥��f���3K��F�W��'9%�{ysr�B+e`����������k��sL����G��4�P���߄\�������/�MWQ�,_��]=ɤ��`��HT����-r��˄��<��-��믯9��5|Rt�F7{������v����Ux e��8��g�'�tT�ݑ
L�t��{S��u��_��^Y*��_+RS�v,������N(Q�D/�N�@K�6��?��kG����4��A/!�w��K}n��ɊB��?�{��cr��W[/.9����ɓj����X z^I0��\a��G�:�f�
�C�����C��G9��H�4C��/��dZ�����w���NPM4�`R���S�,�o3��L1'���A.=��/��f؏�քoe�5׾�R�>���s0+a�_�q1h0ͳ��۠�� ���)�ȋ�5� ��t�t�2�󧩯�ErV���G�ME��խ~s�>:ϙ�g٦@��O��<>�K�+l�$����3���?F�[���+RV��t����4�縦�l��uU�nIMǄ��M���0���#�?Zz)}�,��"�eƗ�7�+%�#�S��"ym'{{ȷ����U�y���]P;�.����>$%�b/��L;��F���`��k�[%���)��S3��팛#��E�޽�f �3?A������ �-��. 2��4���'.nr/���������ƗH�/�{��m��"�Ac��K�,"$�IGƢ��0�Zz*I&���T�_)�Ǔ��_�x��=I#��C0�v+`��]v��G�bA��Aٽ:(Hi<OH�ހ�w�FN���O��AR}Ex"9��$��_�y��Ov���Ҽ�C�_)���_���{�N�Pk5ؒ%�A�����������s,,���4���c��$�H	9�t�xn��w�|�k1\�*o�t�)�y��1�hd���=�mlQ���!FG�Z�R�~�����^NaI�ln-��	���_�_����c%e~� Y$�Ъ��L�������ޡ���Y(�lz�%t_�6�H<��2B��}�]Ҍ�S�����e���� ��0Sz��g�
�&��'N�5L?�[R%.�)��Y/��5����6m�ڒ���Ĝd��p��,!z5�u&���ی���;�h˅Fn۝�P�?�	U�R���~�i��Lg��x�1��_��iz���y��/��)b�����������V!n)>��x��$;�Թ���꫌��>Y�"KS+���2������U����z�)ǃ�v�6��;	c+Юk���r�k�e}�{�������� ��>�xo����	����2`oE>��"ԩ�ۂWj�$$�%C��L�w��<�:���уe�F�8���DC��D��N���ѷ�'o�:D�.Z;��a�/�G��U(����|��O��!ՠ:Ϸ�����i�D_n���a�/?�~�E�P�~��l�E�әn>�u��8�j�0�2ӛ��1��DB�]��e�!/���\����s��Mug���Җ���c(��A`��qF u�����BT����{��?fG΄*�IX��0F��\�+WB53�ɍ�fuy�&j����X��V�Ƈ?�=J1I�4�궐5Md��bn��
CA�� Q��G��Zb�jԩ��Xj�U�Z�g_2�O	��A�b~��_ޯ����C�"$�ڷ� �H<�/4��EcĦ\�*�9�Ät�˦Y���5Έ�_�Lf9n+Zyߒ��h�!�z���RCW��>޴�'r��U�<���ν'�.�~��5�ު,�0���u6�jb"6�:I���î@k���nj�	,���&OD8�����Y^��r7?��m�2?��5M25˝�E:�3!π�=y�O�m����.sK�E~�`0�����Ib��P��f�۵�x`��Q��K,|��z�c���%W����.Lxd(����ڀ�fT��6�����,0Q4�Eqt��x,�A���a�܏|�~V�d�o��a_|t"x��{���n�߀�Ά&D�#a:r�����N�ц}��rsߤ����:Z�JS�� Yd\�����s!:��K�$e�C�׆6����8͢K��˦�������(A�G{��[zS���	֐�*�{Se7:K>����OG�9=���}�}�8�}�;NX8��~���_r�\��`�^&»0ɮد�h�%�X�l�Ҋ�P�e��nZ��>�qx��=>��~��A@\��ߖo����3��դ!�3e|&�&�YY���vѣ%'	���ǘpܼrSGd�h�)�^�VF�i>���p�V'fXF.2o�f��:���1��Ol�c��Pkl�x7O���t1���B�Y��Vz맞���r!휬�&��B]ju.��p-�X�FF<�$6D"R�Wv��H�GsA�J�N ese�Y��JL+1My��-�B��.�Fi ]��� ��us��օ6|�w@��3`����a�o+�|SDp�=��E�wߍ�p���nv�ȋ0A��Jp!��ST��4q���M!)�r&�2++d5��\sf�V���ԭ#x�s7��?���wf̬��('>��f�^�5?E,ӵR�*,�v���g�R 3<_r��I[d�zK��ן�WYqDb��r3�X)�y=�q�<PS�*���E�8+����9�t���������^���|�U�I�� �d��r	��5�K���F�L���u�F��xs�[.�MH!u6
����p zi�D޺l	�阞�Won`(��/��o}-n����Gw�x˧I��8�D����ފ2fh���kk�@>�K��hLn�C��[#���p��4�������ώ}�M)�z�!|	�R�^��(��J[�����������)�t��.�i���01V����̧���>x�u�S�0#]>C�G�=���8��p�3�Ȯʵ�B���c��D�`�ۊ:�����	b�v��n����s�z��Pg�����d���Mѳ��n�h������şc�X��&�Y��H3�аg�Ek���HDE�l3a7�BGh�'L�A���#d��*��.F�vd�5�sM5F����YK���bo�H��=X�Ѱ�)y�(���.s�N�q���eu5�t�W�\����-l�qj�o��y��ű��������� �XC/Ib�O�R^��Pe<(s8X׷�����^^�\�9���L�R
�B;�?�T�Y�ҍ�k��̶}����E%��Z�F����t Һ��,m��!4u��6��Ñ7��{�7�v=����i\��&	\>D@N��R=�፱1������FQkp����TɦA�^W��ۡk�ⷻ	��p��G��ڧ]���������%�?����|�\E�c$?�t���JLbg�6���-@�>��g714��F��Nc ���6Dʄ���^V�&�)G�� z!���+�d��2�lD��Y�Ͼ�c��z
f̕�J�Ԅ"�`��EU�vZ�T4l�L��Ԯ�tA��9?�j�~�C���%���<Ѿ��|�_�%�N8�V(�vK�M�z�Ѽa��wQ�Q@16mV�:S5`V*�Q����υ���O��nu1��~l�̾��y��!K��Ӯ|1�R
�L�5��J�=[q��/u�����|�d�1�[ ���Ӆf�d�C"��%<��W��|�,:������R��x�����D�U|n�vi�D?���n3��Sa�v[X���NJ� ��x!z:��������6�do�+�5��;�S��U2���ۉ��41�E�
�G��O�s�V�v�!���d���l��
_�`�-�A���5����d�V_�~���αc���	�Y�?g:H�\/�%M�°]7޸V�o{�QȒ�{+�*,��.!���Cx�a"�����#	�G��WՌ[BG�ݧ���]�m<�U�j��Z���j@�3g���|��Fɧ�L4�J(|� ���=_�)����t����������4g3O�4!�اEx�_���� q��Q="<��?���7_XT�p����YR�t��Z��c��D~~}-�ފ�iB�&�O���5N� � B'׈2��1�lKё��M���~O'D��u87��,R�c#��z�s_��3��u ?<�?jo8C�f��$#��T�|�I��m���c�J��v��~w�A�!yDUعSV95�["o?��c��q�_�	�Q�eO'yv������Lv�[��^���]�];ٛdv75�N̦�\�a��Bk�d��
�O�o\����9߾��U~<�53{*y��Z�s-J1|v%���8+��W�ߢ����瓵/����A��[����Eқ�j�9�|�COHM-�/���rֽ�j��r�*4���&�o��vt8C��C�։�k�����"�.��D�)���?���#џ\c������Y��AK�����M椱�'p���o��P������i���G��*��U_�Y�o���>KM�l����͏�k��tgB���_$�.`��ώ�L�x��DP�q�,m�
��H�?{g�-���ۮ�� �G%W�FD��-@D��+�����MQ�l4Sp�{$�v��-��ρ���ќ������@4X������p.I�������I��$�UJ��^H���aozƠ3����]�[��~��f�N�sA��4��s�����@�H
/��^I�����Ak�O	���~
��s�8��2����p�e�4��l��q��d��n�e��~N��${%���E1^��_n���r���F�p��f2���r�G��a$6x�׍C��̠�K�'X!��`
�����g�=��hONѭ =o�t�G:�v՘5�d8�H�ك`���'SK���!Me.7ܛ�"L82��'�6�U���DF�)h��}���N��;{��
�V;��D��IB��W�E�D��`ٔ_L�a��H䤨1�Nx�e�Wߕ�el�|$!���!�O� J�gL��R��n�1�ă[;���n��n_V�;�]6��k�fG��?�y \�U<,\�z����G�G�6lEp5��W�����e����rН���7���8p�|��V�5��X�ꏶ>�i\]Ȗ�6S�4H��)�&� v�;񆢑St�e_P��x�ޘ!I�y�CDO�.U���F������݈������ϭ>�f�loɍ����R�����Ӻ0t��dt�Bu8�ȜI`/�X�ցBJqc��Ji;_�%^v==�1��^h5�T�[8�Eh���g������܌�4������	��es�r���%sJ��@!�@���ӝȕ��0W}��q���Z�s-v=3��[Ћ�-����;�J3G#U.��"����Hc�Z���p샒�n2	g�QT��0[��U�v|���W�B\%�m�4Hj�pV���cۥW4�h�+��� A�Ϟ�n�Q�oߋC���A��Z�zn�Ꮋ��X��N���v�H�0>J�r����B��%P1κM8��穳���9�N�&�bҤ�4��mKO>�ŧ����41���v��/"׌�Ʀ������	R�[���/$��Ȱ2����9�3H��8�p;���Sn�12����;!03�I�͒���Ы��������գ��g^e��:�f5���Jj�Px;M|X�k>7�9�ȴ]��cM���bM|@C�u+��r�l��Ik�km���_Qoh,��q%�O�|e���#�n��p+ӣ�Dg{�rV��HT��J�O����D��ү��=��1���ӷ��s�p��RƋ]��ᕸݻ�}��� 77��3�����&	A��Es�3�Ra���+���F*����.��;�[5s�Xa��oJ�!E@t�+j$o񖇻�+-v��1:��ֵ$fޡ�ھ��OY[�=�F�\Κ�N��h0.�C�l�Fcβ�@+ۏ
�[]Vҫ�{�5�uD�2J���uo/:䰨k�c��9~Lh,�3:��;�0׏q�{���\-��J�f�B����/�ٕ@�o#S|�L���"� �p��-u����r�2��yk�v�ҿ����Y���J��A�8�G��g��zI�t������q���7==_'K��]%Ѐ��0��	1�ź1x�B�'��ۭ�|@�olba𬄒c��|��{�h��H�v�*<2�y�[n>��1�L;�֝D��p}�E��W4ٍ�[`#��}�+�����7,�l(ڊ�q5���7��B�f�
�����V�&TZ2a�k�L�8x��?5��K��ٺ��ŉ`��6���'����+x?y���F������"�⫫+���Kj�p���z�aҞ�~�W�̺þ�k�����7�1�y��I��Y�uK�U8�^�j.�z��U�M�s.d������8݅��ꡋB�5>,�3TG`�7>�$-���PU�K�1�D����rm�3�2%�$��������;��w�?�;�ޢivʑD=���~�IZ�A��$���d�ha�yF4�8�����i�A@ekһp53[��#�~����l�W4Axo���G<���7݅�>F�V"P20���r���$
��y9[qV]�6b�ͧs0�MGLܡq]zq�@8v�$�σ��B��C*�����n �g�*i}�~ ӳZ�װzxu�b�gfb���.8�(��qgb�ޮ�r��Rs|ԑ���^�t��ZRv�����j��E��1��ia�9�_�=u�Ȑqӽ�a��Cq�W*���"��l�OfaS!�5;XO�%G#���M(�ENràG����u��G&Z���1��'5�Y�2��ڧ�D�����6Ew2h2�	ثc�
��S]W�|$Y�1Qb|��U1�{ ���H��9_�8��Q� [̎�c㪂)�+x t����[Ȏ�YR��ج�*����g����,]4S�a�!G\ƛw�(� 
����G���?��Y�£7��7��ާC��������*��V��?I�XFIk���z�dXZ�L�/g���
��̕P�E�amC,)ĕ�@v�S���r
��܀((o塠�w��an]}��6yy@�������Ql�&�؀���io�<�͉��/7�-�g�+	����#��'#��Ir+'��Wi;�4�G�����6��_�٬��zj[�S��ccd��?y�|��ԩVGv���1dCb��kmL��pXG�Xj�|\(��GH�(PK�|@(��JVJn��ޫZ7E���	X�2b�l����)eVn6�S&�hߎ�KY@�!�a׺9%R"XOz�GŬ��c������Q�!�/����� S@鳮#�1������y~���`�=��	sQ��6�� Wa#&F~nʇP��ZP<��ԧԙl)軲W//�j=��L���>X`����㦨���RRv�So�	w��z�7�of��(ѓ$�6���=KT�!{$f���/�9�5�i��u�����Ă�����E��2}1*�Y�A�}��m˷.�V��'<���?� �"�M����~#j�����p�1,�H�"i}N���E�tr�i����[WL���#n�.=N��87�*���R�u��^pO�bw(I�@VV�m�}������g�tQ#pRTK;�:��N3��|'�}��Y0�M*�$ԇ�ꥂ"rǃY�$C���}�ƈ[7橥�IZm���C��ql��A�۲7;:�F^��g�
���ꀲ����n1�O�&)o�'�&���8�G(sA��{���E,�t"N�K�pe�`F�΀�6�6�_j	?R�~~����/��ɴv�9���i���l�q-ۛ9'ț9���"@�#Fy�������#,{�vPk�~��]T�㕯A˖��<`����p����8�b�X!��{	��^�xv
2�Z�l��[]��S G$���0)S;�r�R�IH�o�� ��v�٘l�]���oW��w�w/u���m�ql�c*��P�l8Q����L�?"����������P�8P9M�����ś�L�F�(ɭ7�1�H�����d4E�#Y����V�B^���$��ptt���[?��'!a��ՠ��ަo�%Vhz��hjt�Y$�o�&�g�L	��`�����}��{,RH�أᬀ~ϙ��p �lU`��j�Suv��|MY��Zt2��������޶�b�����R���Zϡ_��z��!#�L�R�}�e ������i&��#�.��y�g��N�"��@{Cw.g�^؉*�(��5�Q�5�.�-c��bHw���U���[�M�ݴW�nؤ��*������nh�T���KW�����2���^�fu�f�'��hy��:�㝧��F.p��s8�xb(B�\-�ٖOy�p~n=��[an:�h�V�C%�� ��w��:"�`X&8b`���$֮ Va��в����[��b��2���� �mǚ����/�HUD䋟#^v
\�n�>G�@�����7pȪ�����v\�����aÏ�A�I��G��]�9��$*�y���A5e��/�"�܊u� ��S�P���f�;��������H5�4�����zcn=�z������v���'Cʥ@̜���V6<8��n�_���G��{�����vz}^
Q]��G7n��pR3�"�KT�5&�,�U�i��:Y��� �0R��~��n��O?B����좄��qU:U�J='�V}�X~op�#��Q-aS��{�Az9+D��{����Af8���+V�� ��Q��#�{9��� 7���K���-D���:M��13z	�����D6�/��	�d-}�<*7#_v�G�!T�H54�y��z|Tt�,���%c����<��x��-�
�*\�n�ݗݗV[��3�-X]Z:V��-W3۪n�.,M=K��Us�AmNi���eC�@���[�W��zm��O:����cu�W� ����RU	�{��CK tɈ���޹���A]��ZFs��7���Q4}~���um���X^0�`;���֡�M4��N_�L	�:��~B[�Uh_�`��&�&�P��ۘ��R���x������>��e׃�"�����Y��"�&����ex��i��])%g"������-�Kٻ����y����|��Ln�U.��u�����V��ya�П��E˧��Fk����2u\7v����5r����aP}�?����թ8i�'P�c*�#JPHh��ْ��]�$A��ן�?�Y�>j�u����~�>"v��5�.)Ѯ=���<�B��HjH����C!�5"Ķ���N��~W�C>�ǉ�6�}�v�7�kΡ�uS>�<��b����ߤp}}=933f�ė ��-��=n�a+�%ra�so��:[顿$^uzi��srU��AVP)�>;�B���Ҿ��H7z9�`��5�{]o1�L��kZ}S��s��+���,�t&�����:�R��V�|����� �a:mw�wv�# i���P(r]�_J �P��1�%���<��g��Ӌ�&O[Yn�B!}C,✩��U��
;y��B�l���)�i�F���Q���$��B�ݧ%�n	k�#�hs��^���΄�,�Ã�1ߩ ��vPp}!����B��X|ײ�[����F��l�������´�v�B+�H����#'�����W�g����8�����1喉�( ����K����U<�]
���j��[����d�QELR� �O��u�f����,��kx�)= ���D0sg�2&_����D"P�,j��]��	DK�n�wS+)_�脟P�pE��FւQ��k��m��0�ιg�$a�`��މħ>��A'�u���*��j���@��Q��nm���*jj��Q��XV�g��x�)��S8�~����,�V���}t������(���/��I��0��<��E��**8$�_(=�?|X^��Y>a��04Fʕ���LF�/L��9���+:{��K�4ZL�*��wAx��8ghH�+�l�k��]E�D�{\:D1�JV�����W:�9F;�]��7�8	c��@U�����'�5�76�H��R�����rG}�ɉ֐<7�s��(R����i̷-�������e�/�OS�����gՃ�M2��R�[��)�1�ǹa��sBe��L,�s�0�ժw!8=a%f/Q�B���y�<�=,/�d׻����L�w|��w,b|K��&=�`]/�Ҷ�)�g�
$�?ٯ�4�u���a_9Gޟ�#�9��ޜݫ��^�-�0��ᱠN��mPN�	hu���;7�.�I,\|��`�%KM7�=Y�"�ͭ��E�1����8�2t���?���i��@e���������״��*������=��(�=�4�N5�.?�.44\�6y�՘�3��Էˇ��/�)��{s�Zq5��v����:��L�"���q�G*I�s�)�&������jbl���PZ=�3�O�v��S�{����DYL�
��<x۝�k��M��!* �7O��i��<b�}�3�B�n?)-8�s ������P�[>��맜�Ay*��s2SC��D�{j+Ѩ������!��d��M�_�+��긇ǳY}�c����~~�׌��x��������i�JUSc�9���6��b-"�q־�=L#'RC������^wZm���x�M
���Nc�F�����ew�"�\��a^-�!=����j�S�APQy��~/��\�"�3�?��{�EK�u5zQ��$b��_���Q$��i����� ��������r1��۪ec!�ޜ�Y?ފy�ΔÚ�jf���#!�?dV؟-���f� ��i�ݛ|��IP��3C~gL�Q^x
�h�9��3��c��_`�LE����J�PL,~�����^Y��E���bq;����w�J��@{��w�� �F�<7S�)`j�
Cd�u�Z���j'0���������y�ͧ�x[w�F���#�
i(�p�ϕ��?�cܧ �@T��;^F��?u���	l1)��s%e������y���ض���ضm۶�6�ض��dc۶�$��W���<�T��s�\��LwO�|z�{�
�[�# 0���KrYe�����	��\��� ���ר���hm������ی�%�i���PV/>��^
��	��ң���ؗ�� ��p*"/!'�U:%1�����pi�Ё@2��ዢfV�n��P��e��Đ�-�;0݇u�XF�vKp�Yi
S�����"�"!y����,%���3_���j+	� ���Nt��7l�z7b��(�ϖ�0��]�iv�ӆ�]�����"*�\���@��BK���Na�|�LΣ�(޴ud37������?LIq^v�Q����%Y�����J�>��DCS�Dp��Sr)^LK� �	���$�'�	?A܈�If����#��	�G�"��T� �7y��C!5۬F+�@Q��k��;���ڵןK�~|c�ty5p�i�ط�^M�\�^�F�z��z"�讔�cᓬD����Ƌ���ǉ���!�����s��A�=A`6�4�|P�t���Sߙ@�����5
����,��)^5�T]h���pz�v ���\g���d2�>~�p���릙�7?,�v�c�ʔ��Hd���#��C�B�Ix��bM�6���O?ռ3.��w����Щ:f��r\Y��e�\�3�[-ǐ\H]��Qk�֜���(]�__�IH<toכ+���Q��T�R��	h�hpSe��YX�;������^h����/S��lV���r%����Nϓ��D����,F^�Od/�"Ƹ3��黬ь,WF	�����H���Vja�bp"��E��z��J��DZ�,�Y��wp���&w��L�#3Q���oZ���q��6�Nr�eJ���1(5n�n�ߤes�̶:�a�����z*��\�p�1ή�}X��D�P�\QjX�1��c���ƶԽ[zHCxgj����4�Ѳ�Z���m�p�Z-�3�[1�n�%"���z���h�f���% f�����֞�0w5]��<H�I$4zPe�w�&��b���H����Z0:�a�/ԈÕ�mD&f�8p;��j�1*[v_oWĜ}G \����.,�]���vA1އd+�x*�h�D�A�Rndwy�̍b��\���wV[�[��ۃ�. 6�������I�E.g�$){I�[�.&}�� ���f)qߥ�>3�(v�VM~�@^R��<"L���y�[�Y}`���Q��]����"i�ʚ�זA�ͯȨlQ˩;*��*��%=���h[n/��$�6u]��S�+��	$}Ɛ��p�H-�H��+;c`1�f1�[铸3!ʭ��i�^+^O&<d��5�:Q��h7y��h��D��~���V�v�ek�w-�G����w�ML:@ȃ����y�\��}IE;��P�����>��vF+��Jp?��r�L#x�X�,V#	�}�t�E���(��6�c_��O��\I�HS�Ꙃp��"ꁉ]x*l�_ڐ#R�fť�jl��d��u�!�>��l�BON�KP��I"6����K��h�"�-rŚ%:�p�~���D���3��y5\WˡNr3� !�E��	oFAq;�x(P�l�;r� ����Xˉur8���'i��A߁�����ȧi2�:9Z�h��ݲ�̺&��<�����_�|'�unp-t�w0^b�7�*8�<
7Jvd�nh�Ky��1~Q5j��~��z�����	�'�5iڒ��G��b�#֚��py=�R(��D�t�RJ&�N�re/��UCd��y�ל�_c�V�o������I]��z�&��;�\�Հ7�`9�#8������J�B�|�Zǵ���Mߖ3C�:��V$�I�
�^�[��ӑ��>�V,�������^�uw���v#���1��I��猡y�ҏ��tKM��MMX�s�X2f��Zdw�¾zw&�Xs�{��x7�=Z�"J`	�a�'f���6�Y����"�؉��͔�ɗ�߇�<z�zȨ�׃�	��h6{���8C,�x���V�;Z||���J]���WN�����+�6��N���쥞�зw��@$BVU��Lǀ��B4��ϖh0�M&r
,\T�t��9�{e�>��3ᆦW@�4�]	?��u���i�=��.��~x��@��ͣ;!O�s�K� �w�ML�`#y��G�uU9�U{bUi��Q3�3J��ڨB7�e/�-@l��N�1/[�Œ��Y
�3��T�>djRO�W*}%{&`_;!�t���X6|��R� q`�a3�nKQP��k5���](�@I�B���f�5K��s@rҨ�B�*����Dv�{xfN����CS@12IWk?M��z��i9�x�T��4������D'`/b��[`k�6�> ����qs���e������%�Xh��#+1
I�ܕ��C:�{���C�v���G�_�]��!P_��^�ig��x�Z����n�k<�(�1�z_�ʟ㧁�3AL pȷ�QJ�<��F][6�����1Q����j�&���:V\#��v�̨Ė�o>��:zw߇1,'W��ǌ�ݍ�u���Ԅ��$�ݚ滑�]��Y`	(��@��FHR^��0!ˬ��)�#Ό����q1b24�4���Q7(�r��H�4�7����&�屘����Z0�#Cj��J�W�m�E�<�ܻ�~�Y���T�о�,~���j�I��!�dS��Xɑ�U�'e(������:����|���������R�\���Ɉ��Q�B,8(T��9�K���$<��%&���K/���� �d�U������ͪ���?~&P��>g�F�(ǲ*��Iv�H�&L�ؠ6|E�œ�x��i���Z�mTcA�!��XBIe�_�S��a?-�y��G�Na��`�1�<�'f�&p�CH�4����� �D'(u6v��a+��_}������z�:�W��"ޛ2��:�Yn��s:�:�o���H-����U7QC*��3 �lYeh܉�L�,D*)��p����b��|d�ܬ���x$D��#	�$����r���b�("N2 J��cۥ���PٓZ�i3[8���F�d6�d ��l��J����%p�a�o��D�R ��Mb�X�%���Ρ�Z�w��PL�z#U��G�}�����i30�����RD��ԣ�� M���o�y%��t�X�o|_V���}E+���������>%+7¾K������o��Q'l�F�ȲD���2`�H�]�F*F��B&�GD����?4�k�6�P�R���v��8�?�B�CBѷz�*��ρ�Q�����%	5�,����
3��W�G�wC���n�]	�|��H��������pw{�M���Z8*Kg/���Y���Kȷ�Jo�K���!��O�� ��2B�?�(��=�"������I�맃��[D��~M�w!�p�7���l�������I<�T���h}�}Q��O��_DfS�÷���J��o}�S0�W;5ͷC]������A����Ai4'﫽���økH��5�V�9U���ؘ�`��e�/Ɠ��Fn$G��mq�{���-��wU���[^�����w���l
E\x� �H����e�>\]�B����4C���.�zz��lE�|;����Wp2�� q��=^*
jAȷ�s���"��ΰi��I��l8u�����Ai���O|��z6|����db�h��M[M��I�U>O�Z��k���e̾�l�����E�#R{��[u1�d�Z��s���Np%�uH�ϳ�Eal��t�5 �$�i;S8a�Rl�>�n)&�ш=�C�- !8�*Y^��}L��|�|�I�Jv��~��w&<[�Y?�H�{�07u�,�6O��gc���}��i!,F����dH���}�Z����E=j�.��y�7}w[ā!�Wf�#++;�AN+�U�?@,BpA�W{M��N�A�߷3���>�Hl> `�
�{���x����r9��~��?}I�|s7�7���kypq7�����]�t}�v������� ̑����,�����Y{�hi|�w�䅏��O�A&ya��tX#� "��E
;����+�@���*���:炙,p3� $��&�+��y��%�h��۝2\�Z|Q���79�FC�����Yd�� ���#�=�y��xg^�I�}O֢�Rc�8�҅�i�U��ϕv//�SA/��kn�.�qww|��[�~F|(�iEg0.o����OZ5;������W�}�*��o?����c�p�� ��ȆY�i��r��$�:�P��{=�Yª1wS�p���Ơ k*��>L�>oF$�c������Lٵ�wm|T�kh15P�cʁ��P@�!��D������;�P��ߖS��H7<X?d,�).n�5�F #���e��9EN^��*�B�[�A�+4✂�+<S�]C��ϰa?)���N����?��Ą!��} !�=sLW�����"��Uֳ�v�y������Ɗ���K5^ն�S�K���?�o>���vIm(?��x1���n����w�]Lt~av��G�۲�-�-��EԷ�z� �,��_�ĸQ\����nVD�n��|Ɔ�̵�3�[���ٗ[�t8����ߵ�6�WS�l\���X�L�;(��U/|&��uku���R9���/}�����k`��Y���}�:?���f�\����u����4������NEt�0'����c����Oo%�N�Ӥ��N�nQ�E���T{�����&e�.t"�^Ox�]���J�e��ߚ4
�.Yci���Р�'�#*j<GP �%��<�Ld�A]�q��)�a�p^��iN�^{�U�����_C#>�FϦ�bH#�T������-"�B�(�O ��  �_���#L34i�L�$s��d��;rQ�P����^\!mT��@�_vNAؘDu�LJ]|���K_E��kd���O����AQ%�@�a��	�ճ1�[��BI�y/���"���mG'�H��Fʧs��B[�c�抳�@ *n�+��s�$�Y��3q�&5�N��%�:��������f��M��w�bYi���b9�$�f�jQN��\�����=�eS����ڛi3��*:vRA���XH�J�Y��4�$)���1��=����1�5sz�}�U�����]a�^��6�~���*3����M�9�g����g����AWco�ܪ�>U��+T� i�-W�ڥ���࢒����Ty;�#�<�[����7E[�<��;�V�䤖���Of&&KL���!x���W����Ċ�/�坉a-��p��ߋn���U��C"6b�{�c���=+���Ņ+0{��M��P�(!K^���M�pك<?7� z
��s�4r�z������
94�5n��Zn�M]w�P�<�A���k�}kX��o	$3�Q�����+DN�+:�"9xz�����4
�j"�Hr�#�����Tw+o�;�c��򺅼�7GS) �:Z��)�ss���ڒȀ9:���"ҙ�9R��T�1�<d)}>�4��sT��v���o9�7�X��S��b�F���SGޙp�G}ȥ@>֖�<��+wxi��Y�Q�&[e����p�S�����.ͱ5�y'��]c�j�9�x7��,3(��
��j���wŪz��v�תc�;��au�2�$x7zH�F>[qK1#LXE����E09�'zyo�l<���HL��^>7Օ��0�1�ݾ/y�8="
��.�=m&.ƒ�[�R�|$���w�/{��_"�2G�~�,b������u���H���'CW�!��OS�j��2S/l~-~���{_X�
q�{S����kL��(����!�j/6=��W�{������C:Y�<@�AH)B?����.�b�	6�G����ػ,�����)��WUOS4EVMŔh��� �	���PN�3�m]	����h��+�S%/Qp�j�H���5	t�P�Q�fvQ)�9��Z�4�3!�A�q�����B�p�j'����2�����&�cCWД�Otuח�y��3������
�1x���@B�i,�
�������Uzs8#���#{ofiN�ɫ<��|&C�˧(!N��p@��:O1����KqT�~�(9ҧ<����,�m���1�5��d��] ����@e��ti�G0j�M>�l�?6�0v�d���O�/+}���
r��0^��'K��^8~���I98��Os�o1�R��m�o��]'M��4`N�O���oI�V�Y瀤�-�A�-b@��SB07�j�%ͤAnD#@��̞�"��&M����"�}RU�PV�3��t�q���'�<W�D?���|���~ۙ��Aߗ������-��%����a���5�E$@�1���*�����-TJG�1�U��+'C/.�E7�ʹ�X8�=�\.R??��rF=1�~̑�P�Z"�g�M���˼zmڱ�kST�w�{苂CI� ����������5�mQ�\�+ȏ,f)	�t����;AŴ���Ibt��D���ٿ�8rr����%�R�t��ڰ��`q�b�ћ�(�<�O6�9i��o��H��M���_}ur �q�h��ÈfA��c��x�����X>��
�,�D�	�V���G�Q�6�Ǉ���`��;L�A�-&h�hd햋_*���m�%��m�*Z.C���QP9�I��C�-��(�.w2��;$���I"�>%���t[T��2���,T�(�%��%8U� �VEk_oS����Z�d�k�CgU~��` I�ߓP�ݽVЃ�/��*ڇzL�����w]��GE�GUU�Q8�q �n^�vF®\�.�η�\��w�9fŧ8��)�0oГ�Z;pu9�z�������8�^A�]?{�M0��6��#gj�.x�SJE"P�3S�Q]�A���j���ܫvS���r�ŧl������`���d�Ω%�F�� ���.�[x�ı��|)���.o)����U���3+CR��h7|!�z�C
�a^��iʰ��IHTFף�aW��a�.3Ɨ��L����W����N5~���$��]���b����~���b�L���0���dӿCXU�ԛ��<�w#|cյ�J^��������A���]N2�S���}3AN����f��K�ަK���:C���H���Wb��Ds�L9���At9�v�=\�Dc!S��zQ�o�y4�qYZ.�A�&V?����&h��F�	}e��0�X��z��JY��8�C�tu}���O$u2��/k	�\L���r\}�C]�X�����f�-��x��M�� �.v�*�n�I'eE
k0ܟ���|'�W3�3x���UB)����>���R��2"Ie�$��0�&C�����5[��x0��:�3�MA;��3�,�X	�+�RՋt֗���6�Ǐ�˷�S%�k�1�~��M��ȷ���磶G��{��/�td�<	��]�p��q��,�X����s��(=�,ڼ��5���7ħ��z��i�ʥ����ߑ5����[^�AT���E{�ւI�Ձ+I��_��Ar�I��
����L��E�ѿ~������.�G(�N�*��S���,𸾐�����6�v�Z���"���{If̷H�$N_��%��|�bX���=�
mU�y�U�
x��ήmA��8����}���~E��������q��A�:i _�O�]���s�j]�1r��zy���^���v5P��T�op5�W�s�?J�bX��{���{5ل�CU�򒅠��Ś'H��|f�����_��{k����3�'��g��b�OB�#���Fd�!�n�������N�K�Q7�q��MR�"����,}9|����SH�F�`7y�Q�!��}%@�E��q�m��v)ܝ�o��[<�eo�"?��Ab7k�3��*Y���X[u��TѠ�x��G\qG�F����G]�ӒpE�|���Rz��TE��w�^���P��{�o��A�fr�|���Al�߾�i��z�g�yz��|�z(����=$3���}k�A*?�7��|���Z�0A �sR	+�����S��$����h�_P��#N�rf"�G2�m�F�+��Ϙ&�5����G~����Q���M����Wl�F�i5��t?I�zv�|�bIJ�i�G��c(Y�.�j�q2ﺆ�M��D�o��g��Ro���>�=$�ͦ޴�^�[�b��Un��'H���m̊+Q��*�vqu$��Q���W�pR��f\��K���X [&B~�T��t�d��d��,e�s�q�&n��>K�;.N��bꠄ��y��J�>˲�	(Y&/7i��jY�}A9�`�Jh="�K��� ;�Z�;�Z����ɋu��ܓ��V7��k���㗏��o��/�#���E�ҋ���Ѩ�ò�
|7�G���S[r���`���D���UM���|ߕ^��Ҏy�����Ej�(!��dh�׀ |�����t
��$D��Ѐ�R/s���71���p��{EH��O���Q��t��K���������R���/s�Z%A�BKI�d�ڹ�q���i�[
-��m� ���(D�nǞR�0pc�����d˝S�5���,��^a�Y��x�P�qAe��=�m(�&ltA_��裫�ے�����V�
��tYju��Xx�
�IX�ź�˒.��Bk��P�MM�r��eU`'m�<(��4Dx|��*k���0W���HcMTb���_vd��DټT���jL��aJ��^y�)�p��������g����Q$�B7g��
�_�wKs��D�I��h4�!��4�m=��n��6m��uq���-��g$d�������̉K�)�ItH�߻7mV�UN���Z��|�"�,<��ff������hv�6�ޑ�ao]W<�	|�Xb��eړ|j���a@h�-���Y��ҿ#.b��<P�4h"���=
=�v��%�$x����si�F����#�{��:�ɬ���x��b����#�?���j>>�~�����r�gO���Q�Fɦ#�y0���vȥǢ&�f���IV�bC�X����2�a�i��q=�W���_ȡ��]�\�1y�[+��T��m��u �[�n�}}��B����h��0U�
5�|��I��?;q���ĵ﵈&�򔜎��UC*y~��I_?%�7~2{��OtAB2�X�Qj �vDC	7�%Rj� .����xޮ�^nWi7�{ҹb�6���C����ke���<���s~1��}̛�e����6u�L�^�'	(�t��Yf�m�[L=����`�L�t['�Z\X]�n�4���5�<ӎ�5�(�`L��w͖?1.��
J7�(�ŵ�ټDH���ۗ@�M��Rs*����E��6��W��0�b(���j�(���5틾��$�iz��%�1�[ȫ��*�-����qO�R��-��Q��<XfQ�,����+��[�Z1�[H�ӌ��=�ޯ��tF׊q����[,3��BM�oJ��v�m��l���Ov�S]�֝eȶh\�	�4yS��Y%y��a����!b��t��5\D�~KI'TW�3T�D��2����#`ڒ�+��v݁�3e�E��.ǰ`y`+�Y���Q��ruw��Ӛn�彿����"B����DM�:03saV��^͖�܅4�W<#�s�$��('��O��v�DU�!�����m��KS0i�"��L��_$C0M5-��sS�w���Ǜ�q�<�[�؀N��QﾏQ��+��wnJ��)��T7��Z4v@iv��,�s�U�+ɔ�2���_��-��By��@H��igVs�����h����Y���z�?j?ڟW��?1�$���v%�pE�Ĝn,�l^w�A��u��G�ƒ�U[bϑ����̀�t��l�>&�2�����?�_V�ڧ���B�T�'F�f9�
I���Q�&A���O��;�
*��e�!��XN��H��y�YP-���oQ�>���f"�CF&�eg�!dNU��OF`��qZ%"؏��G�
͍.:і��kF;UNe�.w'����[� %
.l�_��1A�����ͻ�M�(֧U�hB�ۚ�K�0�+vc�y��-�������7�V����SLef��䌅�{Ad���% �B��u�{7����-���dS1H^��u�Wp�u�q����V���/pB#+z���	�)�*��gF�; &E�_�.׉۴�F@�׾4.*�!�s���+ά*��m�k��R8�[�Ex���ti����̄�$uLA¯#��)0�TݙF)�bID���*eN�)ص�^H6��1J9��(REw�O=fSt=�1�-�Z�rZ�ba�\ixZ.���p�X�cT��(]����D�}'�hS6���`oc�!�E_�c];hT�/��Ha��fq}3a�� |X!�ݸQ[�����q�(y2k�>X��9�X�m?�H9i��w	Q��앷a�R�O���*�����Fʜ���g��7��yAZP���E��bb̓�6�����Ii�ۍ�G���w�OƝU�e>n�	���˲���am�xwr��>���c
{����N�ޯ/	��-E)4U��Aw���6����`h�0=�d|�JL)��_@?}%H	q䇓Cv5����lN�h;(�;���=�L���a�cG���qh5"�'1\���p{U��b�t��
�[Y�b�r>=C*�'g�?�^�j��n�蛵|F��Ct����Dc�����-įU�7����va����I�hr���(n�c�*��K���N���4�z]姙�i����2kn6�u��)�R/�q$wOOpɎw忮0��Xx�nnq�٤�SB�^A���v�X�8��V�V�1��T��h��B�����O����l�j�y�s�*��)�N�7wI�Ri���\�!RR@�N_wz� N�E���{�[1�����������N��U��6�)��M�8D4�2��,č����4n�$C�́�7t,�de�S�W@B}=>e*&�7֜��I0�,�n��O([n��f�Ȋ�]Xv)[��*.�v(���k�'rjϸ��zv����ŵ� ��4R8I�7���`+�&�c���Y?��r``Xe/�^����ǥ�F�sl�d&똧�rce���b���r�jqGiҺ��K@�$�:��W�d��Z��}wuQ,�c���h&,K� 3C��V)��F?�*�n���&��v�R��sG4��=���r��=��=1X��c��,&ߵ��J/���tԨ2_M�*؇Ǚ�	{x����ȝ"}��j�8z��+r�R���`�Q�p���+� %%�\��4VL�)�Η�k$Sh���N���_ˮ��߿��q��a�h��-�(%�@1K%d{����w����Q9af��z�:���g@��щGW����6U�T�:u��<�-�%�\�X���;�}���%2�HyE1���i�O�o��lNG��uKe��&ay�=c8���ª�+���U�l�G����M�`ÎF��_JA7�UuTW9IS^����w���a8{������̭���c��3�P(��W��hx��Ag[+�r�.�K:�������� Dөx�?x��#N��<�l-K��$�="��Q������B)�g�=A��7����$����2�n?�3w/�[د��i��G\P���\���>�\��*��$2!Tl��(��73�3�עL3�I��$��ne���Ryjg���2=s���u�����G�<!�k�����V�\G!nm���� ���N���އE�L��⩪<[ �\�Ɨ��e}�����4�-�DN̤����-U�.�s9"�`P�2&�����z8���IsIՊ�V� ���^�E��K�6�P��A��h]��B8�"��CU����u��i>}��Ƴ�����4�Ѿ��b�����y��x�=vS���F7��;[N)y���E���]�0%�>�=E�v�4�7�o�7�C���p�y3��`S4�HM���G��hlx�xA�6q����zk��d�-P�؈��N��F�Gʜ̤m�9���l�"G��R��TQ�i�vsI&�U��{+�k<��}�i����޳Ηx�p$��v���+��6-
%EJ�9�5��]�g�о@,���x�3���������Q��j^(��� ��B̸�fp寵��*lIFL"�S��r��3
��
veh��{_+�K�F��帞h#��1;���{���ƙ�*z��5�%;8T����N�^ �(J��i*Ӏ�<�.9�Ȱ뉝r@ ��2PE'�q������bE�I�������)F�W��	2��t����i��V�� q2�|ը�|�����c����ԟ�Nt��h�x�����N:���7���q]*޿{��i>UL�NT5g��ҁ���Oك���u)=0_+MuQAI��9��V��?6D;�ӧ�DL(K\%��_ӛ����ո���X�	�B���ʾ����J��oS�d&/[/�0@"b�ӕDpz-5\�f�f��E�/.vG�H��mP�9�����O<q�iuݲ�)z��̣�V|z�A���q�kݴ�?�р�=���m�j���bz7܏S#>ѽ���n�$u����F�N�f���4jh:��ܯ������Q��3f�ܐ������m2Z���!�A�j$D�pzڈ*���ԅ���`�!�ӹ�j��jPsE�?Q������)lD���X��k~�@���b���飵P�Ѝ��Ș����*�RM|b%;�	h,��[}���ُ~6n�]N�n���m(�![5�E룡�bVc���oRGK���"�ŋ
l�ՏN���ߦV^�z��o�Y�?��V8g�&s��ސʑ��Ҡ���[����Σ�b��+/����2��ϜaȾ�F��Þ?Ѐs'ќ���,�]�d�%��R5�ț>g�	0��a�](R�c�J&��=�oH�h���qzW��$�J�=�L?������2�#�Q�K}��V�n�e��}}Dk�� ��e5rq ��e�z�n���^��D�*!���	(����,���2G��ӧ˸\�:���jዳu,�.���(Q}����ˀ�Oس*ICбn�6��}����/^9�!V��|=n�C��Y�CGf�G�"��ux)��!P^c�	{�l�~��RJ�X �k_NO��p����3L*���E��K���:0���CX�h����L1D���b��)m��`o7L4E4�y@��d�F9���V������Ў������8���rmV
��hp8'��Ҷ��j����5u�v~Vܟ<v9��VC11���g�F����9YmrOFM�9�󵩫σA=�"H!v���fF��CE�#�x<�|��g,�P812��l�4=ʚ��&�o��W��e�ǫ'��-�P��K�-�����?��5d�޼�pgt(�#э�Ő��	�4��6�a���1�rCMHG"�����]���V_� �_�����z>`�<���-����E��e�TNgP����%��	�%�O�n��ԉ�G*��k�{YK�
�;��6�dZ�pC�n{*z)B�C*^�eU%��p4~�k�)*�mj}{���~�k�1V6,�+�YL"@x�|�C$ SXӉ.�<�P2�_ b����Z]�s���ٞQc��������r�N�� �]��X������ey���A��=����փ�Ǹ��ceO��)� ax�o��'|�]�戤�j����`�G���I�u�&�=8J���F���!f2�%y�?ܥO8Ov���xu��"Hy�M�b�<?�ע���ɤ$�^�BՄ�	iG�ƛ�6���O|�!@�jW]�+����]$�_�_���$�%_7�PǑp�UH"(<s�^��<���-�6��)�e���	o�A$u�3��-�\��p$xv�-��C�4�~��x{ĕh&���u��D� �*5%�y��8��ȣ��e��M�4Q�݊l_�����w�˚8$�64?ب���k�t�Ѻ��Zr�s��b��ꨏ@��\�}�~����\�[��3��a���$���v���Lǚ�7@a5U��[�[�Dr�J���i�ߞ3���yY5 1�`^G��y�|py.F� �^��[�4/=sOV�f[]-~vI�ƞK�B^�П.k�(��[D_�!sc�i��ݜQ��
������|��_j�C��w+�@�γ+�i�>����E@��z�BD��f��w���.�=��4�ܐ���w���gN�*0���j���D�A|̹g܀(G��{?�JŶI�2���j~,[��]/^��5~�~qh�N�J�}���	Ȉ�,��&n�H${�/��JX�Uj�@���5�w�2+RSV�s���$.PҢ;]�'�mDR(V��_R���us�|�}er�uz��b6��.�%��#êipU�!D��w�z`��f��i���{��@#bs3���I?������+�F�*�p)5/*��.o�<��U��X��d<�� �i��7��ȏ)yr��N�9�6���#!I���n�S���;_��J�'��gz��&��?��Q?�[�����l�H�5t�N&§����r���e�Ӂ�3�}.n_W.�y��!�N9N�
�<�o�ϖaS�ק�3G"����F�����k�jL�������0P��mr)� <�,��x���9E�
��Hp�Œ�U3x�2s��������$������	�o��j��2MqL19"F�%k���C皢�5�v�9�m�Q�%[!��4A�r*{��@�`j����>N�~��S�ޙBƀ?����6��0"�_p�������5�y�L�U��2ߌ�^?{��5�Mbg��Өվ��{���u@���]���ֵm�<_O	M_�}�Y����irM@�(��Ѣ��oa���/�;��C8�R߿!�o�;���K�h�5�Ԥb���7������1ڸC+��H/��~NTi����~�l{�khg��K��^d��	��ˋX<�g����G�����.�[��l����
���9A�����2�O�V�����-P��쬙j{����~&T�Z�A���9�K�[JT�^)@eG�`� ����w3�w��Ĝ?�k0Ҏ���:%A�ݟ��	Z�"������^�!u�v45?<*Tq������ʺ�}ɉ7��ZD"�y��X�t�'O���.�4p���2�(�'��6�9��	8��E૭
u�U��@����PT��d\��dqG�ͽh؄M��+�@h~�Pq�F��ph8�R,W�k3�,!xrH�|ڂ"<�瑑� �� ������ t^{�C'/;ڸ���������=u�@�f�N���k$|,j-���P6�ym���>��
�h���:����7a�S��*�u{ⱆ����{u_���� 9�>S7�)k��0vJ��1n*���>6�/�ք�Hs�t`��5�XPY�k�V�S	�[����w��W���i.��PX�A��G�->8�p�%Я�����)i��q�Y� B��׋[��l��x�pGVg��//����;�+#�(��a];��S[�����8�nA�iHr�B��t?,s�A&�d��O�E�����e����p)�R���ƇHp�<{���)p<�2��ݮ�Od��(�V��݂���^�.^O����U�i�H��G��O���U<�v����Z�'�Hص��TUE���h��.�����4tgϓU��}�!��X�ƛMȢ���&�"������S��kC8ȗ<��;$���>����d���2h��tM;N,��e�ё�B��#�����ՁA�##���Z/�+��<�y���N���6���wQ�y�O���-�>�kt���>�:��`A@�����@I����И^�/K���.��k͗��$��.&ܱCӅ �ϧm��Gk�9EU�Xw��.׭fG��~�sX���`t6[�w�ZQxrA9����ޥy�or��_�����(���Ȩ�J�!"g���������;�e!%�{�	�r��Z�����k�@[1QO�/�%-���M��X곞]TK��RS���ؓ7A������:Ɖ[�ec[Tg��r2��.��R�B��qb���`�C�f6��nm�!]�}�@��Ҫ6f�gS�u\����EP�����j���;�FY�ã�C��D$66��3J������t,�x�'�����co���s'�7�����ai��'W+F]����-�oJ=>��[��^Sa�v���?����`�G���e�����:��h.k�5�n�dMKR�HV�(
p;|ȑm��T���AV��"���C��6��3-R�".�H} `L�PP�f0�
��"��R<�
[����O��f�2�8�/����.[�,VQa%�@�����Eph��KX�O�޴�������a�3i�el۶m;�ضm۶͍m�����ضO��qr�w��QUOW5.<A�v��@@w���W���_:7&�1�"�VjRdhʗ4s����ט�T�j��O��u����K8Ë�P��^�x�u�FH+���lY�� �8ד�MMf��x��w�:nU��Jm��@z�2��0Lc��g�� غuw
�}�3����J$7����區�YqE���p`�T�	�ۢM�KNC;0��Ậ���</_K��'�y}h2��@��l�] xhDA6���*��CJ��wHDH���`Ԫ��VԢ�>�"��5�N�]7.�W�vtk*�����̪*��م����b�����_����k�N���n<=��|�m�jC&J��W��yܴ	��e.t�b�\X]Я5�*U��U��xdp���jm��S+��m h.�Tf��
�k�A��IX!�LCM�e��	����
��Pq �9���>Wqώޅ�H��"X����!#���`�<W�ё����&CHڅG���6�d1#�7U�B�#����-Al����kq�݃��{	�큩,�����![M���~����F?����*4���ti�@"v�z}r���Q��~H0T���>��ajɢ���t۫dSR��ԡ�@���wO�~N��w�Y��E��?���F<�71	 в���=�a�SR"��,I<���봶��'��"�B���dK��9�Ý˪�h�j����E�@&�e�*��x�43>@!tŎ��a�Gb��Z. �^�~J2Ӻ{GJ��,��Zy]z���������\�xT[@����k��*��.�ip�@ �4/��|Qk��zw[9��+��u��Q8z6<h�U���f�dP3x� E
2�
,��cL��{Ug�,�RB��+����1��>��?I�3T��=�u�zJ9ϵg����=��i
���6�4K�ï"��a�L�4^����'Z�*�"�{o�?�=}hX
�����Ԩ�#���$�|%#��]k/�����kt�Gnw��1�˥S�55Zb(h�2���q1��r��N�����H��>�0����"\!���	Q�Gm�1$8fv�e����������#kw�_��]��\����j��n
��x�dz�i����.�w��(Z�S����y�&�A��/��@�Z ��'����q�9�!_�&)�"��M7V�e#-1Vԟ����@����0�^�Z�!�|o�Zu�;���j
-
:� )3uC�Pe�NN����	~U6�7p���׃�+�Z�����-Mȑڤ�1�����g3��Ϥđ��t�?;��@_46)v������:u�~�\	TT ��xDP�ˀb����)*h �)�J���>>������:��\�@�����V��U̘��Sx3[ɖG>�ɦ>㤠�/��#�bӘ�l��ZID�û�1==:�@n�]Puv����ڥ�A�N�ֶM��ܖ�h`;���`we?���2��H�����dؐ����~���W��yx�m�9{2����kFe☛�V-Uǔ�Hzg�knk����:�VtB|5���{���.�F�ʾ�I�5m@ 65�YI�Ή�D��y��@ ��|E 2E[m-�)��0F��˴��v@����X�%��R�)Pޔ�����L����-�H|rJ"�;N&���nY�e�,�N��7��������S7ޥA}�>W�%P�`�t����8g֖n~�Y�Um̂'NJ�}#�J.iW� 'rv�ς[Id{^Bl"dȴT�He~�.& B1P��e0=.�jo������
�s�<j������e�&��Q�t�u��1/_�w�Q������GId����K�c�����܀���b��)����!'F��޶�?���$;��V���Jmo�g6�j�qҟJ�BI�8�<I)��ǡ�u>�S�Z�~�H~>A};0��aNMf��u�黟Mc;O�����#;�L\n.G:R_�Ň_*�J,����fҨ&;���q�a��`mnh���6'&�����oA�Y�-P)�.¨m6e����ܾ�t�hP�0���î<�^���u��1�ޖܽ��xWl�NXeD�g���J�h�qsi�郏����L�Mc^!�m����X�_$l�)�յKs�EVe5�����ix���7�=�/y��kY����>YN��]�Gﯦӯ��O�k���Ӿ�7�D�^\"1�� ��_�A`Q�T9��L]+>��\�����T��E��WvSf��H����R��ZjW��?�[x�34�Gy�4V�w�|{*�q"�� ]h@T@����)���y���PAe|^)��<.�+B�C��ߛ��
|�_�5���x��Z�bU����N����9�*q��R�]85��D�in쇵����+a���#s��A�R�f�Z��0�����,�|�a�h!=�~g�%"�C�����נ��]��Pf~U�J���o	T�s&K5upVg���Fw���_�l�]�#8b ��R��'�^��K�7��^a�wd?�-xr�c�4,�Z�7�B��#��˓�6]5�M�����{@{��,)������EY��]��n���t%�O]2��R�alb�)����j�1���I�Y��l&���*ܒBh��lQ�ru��Mw_��:_�q~�2���|�g]Իfngڒ,��^�ۣv�N�,�gBu��+���i�9Sw>Y|���5�!ojȆU��ऊ&�pP�<���߰{���:e�RǜCB�<Hm#X1b�R�����S�`����G8�i7`z�
���NhN(�#����L�I=�/���Ǒ���=�w�Z����'�x^N?��'{5��w^�?*7S���Fc����u�{��Z��iM�/aL�(Oȉ�#j��)xyє:c�ub#4���E,F���?n
ʺP�|2��1t�a��cy��
 ����`��TA���BU%���Y�ͮ���Qg���G�$9H
Qi�`�y�"X��j���%�jU][�_x��R�M>ݴ������m��(֞ɔ�:gC��5���j�`�nK�b�s����iI�Xo��D���̂TǬ���~�MX�L���Y���B>]T�f���!���՚5��F�����(k.�����}�v���V�?L*k����k�9RYC�W�Ky �o^�"]��O\�
Y�e'���tŭ�zb��h��x̑6؆��C��`$L��@�N7`�f&C���p��E���0�s�`5�q�"�@�Sn:���#t��j6ӶćL���Ó&VJ��S#U�<��p����*(��y7�~��r�L`N��Es��o{+`�4\�tw��Y��G-��vDRd���k����i���5��/�t����&أ:|ӥ�r�y'�{����ПY'��?:�L�� n��0�A%������<�o_C��Dp"`�;��'��l 	��/����	u��^u=�8�J=Z;?{��4{rJ!���h8�4�5OΘy1r&���ւ��|{W[�q7tTx��Z'� m9��߯>��th�l^���	GT~/��� @��YYQG�u���o�m{�J{C�B�Qi���1}���䌃�|�+��R[�=|��'�TI���55�8zR��D>�񎒳j(t���k�Y�'�Tt�s�Hs���������F����&1֒�����8!��m��!;�/�iY"�?%�^F�	��O���IcZ&<5�������MG��A��k��ࣖ*�o��g8�拄n(o:*����7A� ���$�n.~��޲S��g�+�ȃ�mk�!F1�s#���m~m�w��pvE���S<�NJ8���,���2�5G)$,�pW�usB�(NH2��u������yM��Au*�h��U���j�	3A��O�S-��u������d����4� ��Ӝ��K����r
��Џ��(�S� o�*��g �۸P���u1/��?ONV��DϤ�u�E6�[��3��B��fC����Б����'�����!I+���if�13h[霅�b�1�O�(�N[:k����J��ĀF�
�[����0��E��D?��D��cv�k!b�H����`C���E�BD���F}E��8班�:��~�*j��*l�i���M����Ci�	 �4Ј%��AV0V�?��cܞ5&Sԗ^���%���z�Ƨ�F�A����3�$�B��L�� 䖁ǻ� V��O ���Y��8��x�)wmz���<�Ln4|��m���Aq��0.������C�g��Z���$
�,�	��}����O��--�*��D��8����%.��+i�u4���|V�;��f��iɆ�R
�HپS���\C�x�$�#7�-���?�:	Z*?�T�1��zxCڰU������&�x����z�,H�|��#`��k߱r.��4����+�qI�����8�CGʅL���l��&d�T����am\������0������2=�ʳC��WM
MҜ����v��;s��l@���w��p��J����*���2-gQP�HK�>��Ү*�M�S)��xr�hf��&� ��ݣ.:�8*?z�4L��@O�u$%O�fR*��nڌ�}%1��d-'i<2Ĥc���u��
�x�������N�!�6�F��n���ނ���M7)����żu&�K�^�nq)@��V��1����ʉ�<\q�E�!��C���vi��q����Z�DF�9���uS&W	$@d]=��������S�|,]V�gCf�Ƿv��?�>.��.�E-o��0��y�P��!�Z�c��T��Ѧ�2��	 $���ȧu���$)�d�2���մɠ"�UR�%��?�YN�s0|�y�v���RT����˪��M`�Y|,�G"g�뤐q[S8����i֦[��&�(
��7��_��&�ח6C,4y�.�h�����m3.�G߮q̩g�r-Hx�S�����Z&���n��(�Bf�*�-@�	f赵/�k��/���R�']�@�ѩ������{ھl>]��k�4���=!?��|0u̬��Oo����-��m;e�MF����z��	��ߜP�o��H�U�r���ȡAM%<�
"�]�q�_ki�H���$%q���
q�]1�|Y}��>���Fp��0�v��-�aO���No#`!���a�k�~����k~,�H1���9���)�z���Z��e!����/�$��uuweP
�����6���3�����3$ ����5E3R�L%��t	��FN��ɠ�ٸ�"������M��!��'���r�3M�� Nb�Y¤ض�?����0�Q�(���K�p-#ASzϋ5\��ߨ<�|I���j�J=�=����H����[��r�v<^���m�z����9B�9,��R�٘>J�A�f���jT�GSү ���`H���:%l|px�p�ԩ�(�-n�F��3}\�-� �9����Gr�J���a!�2?}VЊ=Ԁ��6&¢m)��0�%Q�<T��.=ֹw!V[Y��0����Ħ��I݀:v���ãaK� w���	d.�bz8'IQ���G?lU-�� &��{ا�\U�k�d��5nC��(��q�g��0�e��2��[L�{.������/��;I�{� �x'�benK�1'e�#�S{T���_�Y����ڝ���6KB�|LA���#)��I=���N�Rn��`�����'�,Ψ�cIq��V������{���8��@� �b�Ĉ���ϙ�粳��.5������	�)S�Þ��ٚ2 P<ya* g��P�N��P�'@w�9����~�,���!��5���Q�Lp*��d��R�	���h�?��l��*_cg�)jeY��5˸�ui^���%�LUd�D '�Lź���3�h C�|�P?�:��E��6����BIp3ư�䳻L2X�8�SM2IM�R<$Q�6��E8��#������(��;k��n=:���k+��nD����Un&�VMDrݘ؁�]������k��p�"w��n�����oO�6d������_՟���siG��D<g�k�өN���1_l�(0�|���!�S��&�����'¨�h[�PeK��*	/�D�u����3hD[|�B	y��B������b��)����N_1��[w��R���(���`Ч�l����V��S*4|��t��g�+�B���,�2G>�7[p�KK��-�b��v��ڃN���50��!���ȵ|��e$�`��ć{
�Oo>��_-���;m�5��Ez5�@"9���2���!�2d�!��fs�%�{���ۋk����l�b�;�jn"� ��?��O��fw��4?�|I�fD���HY& D��6aX�f�*U� ���ٳ
��k�rT.����S�/��8+���=X��}�t�*r�X-����TV��eO�r[�<ˏOO���緑Q��5	�iE.��\�یpgT��Ӌ:j1���G�K+����NT^Y��܏�g�n��Q��w��E&a�_�d�F�(��GӨ6�u���>}_d�-�o�@�6�J��D{P��8����� �
�W��'����>�V`�O��<q����#j	d�!���\�{@u������e�l��z�����6��	>iL��e��Y= *�s�������N�m�钀`������j�/v���$��FQB��fN�`n��e�duygJ�{(;����h�fޏt{��2.����_$���jΠ|��x�����Hf(�kǼe<�S��9��s��a��Fd�VΑ�� iӡ�ح�*HR��"�|�Л��y���`qꜹ{�H��ZCm���߂�?�v���a�������ry�#ď��%�W�9���9���~�m{�#t] HftE�4o,ԯ����o�~<o�|���~��3_��r���(Fw�I�2��q��	 ���d�B�3�f���y���y�NR���fse�]򋲺��q���;�_W����H?�h"�05h!���������Ǽ�
}�����˺�Aj�q�Xc�>ׅfhqu)�f����R��_�\�2�x��b?y���,Ӵ�u�!Ad$�4�����]lP��*h�0|�>��t+w���l�>^uf�R��=��J��A4dL���T���R��5�����vh�³�+ī*�m2e�V�$]�Ic	�q�a6W�cA�^I���n^�yM�!�� z��r�< �_��<���1~c��%l��!�"�W�?������(Nq��g�v2z�]|2���ʀ�G^XNv���w�����~��h����=H��{�-� �W(�x�^�ۗ�b4J,�w�H&6�-��Քғf7��J�@ ��4�#H⛭�>%%`������x���`J|n��+�+B���^��۞sO�W���$�ݬ�'1ށ((���NY=N�ɰc~��
e���#�{yDL�9�,iq���E~����}��`��l�&����4:�0�R�(DK��g~#:e�����p�ԫ8��E��?����4$������g���#DzMX�a���`���_��d� j�� ����lY?�C���>~]��-��t�k�<]#�:���E��7B_���B܅;��l�'�~��9��C����2W��t��N��@�}�-�"���Ϝ
�O�P �6�@5I��q� �=�α�OE���ս|TZ���(��s�>[�9*L������tE�B�#��B��� ���H�%fO#\�%��֦ک�a@�1� �I��A4���aF5���c&�L<�>���{��?]�N$gB�6� X)����]�B�5z,���t�v^�*GÀ�LRD�6�Q����;��Y�"�X $���#�c�� �+�?J�T"�|�_��_ܘ�f�>}���-�-͢��ҍ�����Hnϖ�$d���O�E��O�i�Wj�MǥV9y~��FZ(N'�'����S%d�pN�<E�R|��y���љ�f�S�_r�[�%�*��*TC4�&���
œ��
���v�5ɭ|ۅ���Z�td(Wirp����q4_
�A��c�ǘ�%a��ƶr�>Utl�|
�_���i+�?�9��&�g���D��%~���W�j>�Btφ�s�S����&�2���s���D����r;�4b�͉A�.K�x��Y��+,N��v��ϵ����E�k�#�$~B"��������'Q���n��2:�_�V�s�A��P�`��2E���M_T+�1K�����9yep�:�J���4k'�\��,�E���Y��eX�����:*�>H*Je�'7k[��X_�K�vR[��۶C���L	O���ɷ)�f���Qz��ѕ&�ʄ�Y�ҫX�� �A��=��4����'��6��Q�d��S�O���LQ�8<�z¯}��P�=`��lF�ˣ[+��U�o�!�"��^��������T3���C�����^�nEj����J&y�L���v`Ѫ�%�X�P}i�$�Df���pq�;y��ٕ�F�xJZ�;w�b8I{���Ł��d�>�_p�"A�U�Cҟ�8%���V��<9LK&8��JWή�H�n�S���H(�����"q>�q�L��a��@]�Ƭ�#���-��5ax��	�9�W�7�X��p&?��_��e�\1@o�����{�#j��.~�t�K�{�Kl'���7��`-nm{�9��_�%�n�ߨn�������ٌ(5��1��&��p!���R-uW'����M����o;��j;fF���"��Lp	K)hT��@�a/��(� �puS����1���j�Y���N�O߈f����'����vfaa�+9~���Mf@�x� �/ FXNH���``�}�ClD��x�'�{��T�8�GGe^���T`b��q��+}�����m��Q��B�U��xM�Zc�u�\Tkl���Rhd����o���R��ɦ{e.|�����B��׬P��7+�~U�@W�͑�O:��C�
~�q"�K5~̓ΐ�l��0z_�_&��/.�Q�!~tiU�-;��_ �F��ĳ�z�t�}��"��y_�f	E�˔�i�w�K��ݢ*<��8x�ٞ�i�_yP�/�Ȩ�L���gd��!��X�Xg��&g	�a����|�� ��QȌyb���/�AR��ǻ��T{�# ���@k�x�w�*����&��������}���y1�T�/p��⬣l��H�#Ҧ઀Y.�cD��������W�V�A�x�%l��RE:��~L�Ya�}��U�=s���9|$����� 5�&g��H󲂂o��/�b�a�ϕ%���}��H�����- ��~'����*LF��������6f�����h�h~>s�I�sϓnX����,�#'[cVΪ��}�����+A�:}o'��N	t���z��nik�Te{��g��x���Yk(�Ɗ�)�Q�M�Q/w�tp���k/�J5�%a/�/n�'��d=\>j���Y��띠b%X��T���p��I)JljA<֎��Y�8���l�e7�l��qGH�H"�|���-5�7�!fe5	�5��/ءi�����A�t����o�;�7q����͟�����S�j|^Th������L ��\���-��K�x�9�OUq[���oq[Z�	�"���ߩklЦ�_:�����C��R����9�Ju}O��;�JMl�%������pVvk���Th/�U��f�UG���
�&�n�� �,��@M�:J����"k*��e�,�E`o�X����S��:��'����eT�����m˼���u��mݷ�Ղ�G}8#]���1h{���C�>~!�B[��x�E"m�%>[llt�]=��S��@p�W��ϗb̐B����G�F���1l!�S�A�aX`�H"��M2��?m=J��º}�����/n���='/�r0�V$�#oq(0��r,$i��LGlE#������.q���=����F>��,6�0f?�ѮF2�Gĺs�&�?3߱�&��D\Mـ�1��V�.R���T�C�,�B�H�ڇS����u��R	=7�*��$2'�W�X�9���D	`�hD���M���������5U��"A���:dL<���Z�z]/���JMI���
k[���9����� $ݝ� �|p�"dQ���P4[{o�7U�Tx�f�N ~A���)�L�{ݖy^�y�BW�K��Ft����=�� ��FXGlk?�b�Z��K�A���Y?n����������Y�;�c�go!�$�)���Jja�wD���X�������+����b��&1�����t�U���.~�bR3��ʔ7�\3<ɢ���ɞ-�r��kT�y��Ǭ�w��az��d�"����]yy�7v����b��۽��K`�Dz��f�Bc}��v�*���.�p'_XL@!�&a�k���"ؓ���FR�7E��t��G��ѶѶ`!ߟc����n>AY[G�LMG�%�`����j�2�u��G�[�N����� ��E�y��"hd"��WV�ES�f�肩h|=⡅,=��d]M��>W�l��e����X����қ��)�"��C$��	&X��b�t�D}�oB.��z���L��݀6���UBF:��^ay/��|$B�咃��K!�[�l��:�Z�W�dQaRB|vXۀ4L�tV��T��	��P1"��IYeGx扡d�����Vl-y����X8��C;@W8ҘrƩA����+�NbjJ���#8��[֌�^l昡v�;�O�)T��3���x������@_j�=��uv�7�J�Yi.�	���PC����Gg�ln�H<X�yoSР=3cb�%��lY�N��2�A!��>J�����#4ܚ1��T�RH|����lra%���O�7������m�TN���ח� ]:�j�$$�~?IF!�%ò�KZkw,��V	H�f�7#�6z���<�|3�����	y�	���bP�DQ�ۮ{�L�AW��l�Q\�b������n�5I������{��� �5��X.Ŗ�i�}>�蹛�]VU��mf�8���ה�q�"����07Ŋf~�6O��+q�;{�{z&��">�)�=Qv��ȓك�C$�??��4�R�MHO�c�`��&"Fj�ЧE�^����B آL�8.¢�g�,��^3oCO��軒L� N�| ��`ы�nʙU��K�脭�g.����P�J ƖW�)|Z��Aԋ�r��<�4萣�-	%�~�_C����~��ȧp����m���鷗ws)���ZRy�ߞ�����U�3,��tYݷe��a��/M���*��eT�f`x��H�y��/�f�uè���*�َ�4���2̈́�q��z�E�\w�gd�s�2�lԭ-�Z)ܱk���5pU���f���t����5�~ǣ;R"a`C*��qb��v��W���p�*���k1�Vo.���1�5�U��9�DTfo��9���A�kU���kmhQ%[����ӾR㑱?{lj�j`5�u���e<ݑk�|��/bk�_e�ɋ�7a!�}�K�9���	!բ$C��kz������
E�x�����\���?���Rׂ�3l��
z�S����d�wК��T]l��߱��(ÆC/Emu��O��^q�2�0{�
�FM��:�܂rv�j��=8 ���G͠�;�I�Z�Z���

��_Cj�{�w/�?s:��w��k�J���p��VO�Pl�TL��+k^��c������\���F|�ê3^�]n�'�_J�⢇�i'�	�[;�?(^�.vܹ��0<̠�į�
�)>у;h��~��t�}�6���ףġw�6NG�  Z���lQ~���V�.!��fr|<؞	�CW��s8��8�~
FB/�]?,�g�pa�r��0����Vt���
/�}a�;�W��U-K����;8��w���?�#��:�qP͇��dZO�)��nM^�^ك��nllA%\���t�P/���;�֕�oZD?.
?�H�2��Y��Ȩ^HKg5/��.����H����`�׽ɞ=�y�,R���l��ag֕�b}�pN��j���d�n*�'���iS�����W缹�޷��:y�?�c(H4�I����ge��E؏���r��K~�#�IקةD̦G|O�����˛\�x��^�Z�n����&F6�$%1�evj�¦[���Cq5�Q��p������x�\�z^�����",m�d�P=9�+��V�4"�+5/u4��&��O15? �$�� ����G�����c/�G����DW��� #�%�Җ����ӢѼ��ް�jb��X���6aOc& ���K��~&dd�����v��4�b[�+l��qX�X��0�g� �nm6i����J�e~v��00��ز�E��������P<�a5�0u�r����K8r�x���H#�����s�,�JJ>�	�|/�U�ʚ��*Fոo\v`����s��z&�R�#L�����+|w�S �Ƴrâ؇�S�e)i#�s���q��u�.�ϻb�o�1����_�y���@%b�ҞA�3� �b`R���;J��A  ��8xz/Q��W[��j��h��S����Ui!�6��ruv Ը��
�/�����uV��������UB�*A��`ԭ�/i��z�㫕:_�(�4(�$�"U2�
u����VkЪ�*���<�7�⦋+]�Jr��X���bt	��X�-
�K�����ɉ%�H����T���cG�5\U�潊���'\ -�1�ϯ*׬�s1���ڋ[_�s�3,�h�=S,a�
ĳK����1����F�uMFg�O�?; �8���	� �p$&��R7h���Fd�~Qn܉��讶�\4g8���zU	j�G�Ea��NK֚x����i��#}
[��[P����G�x	�kB����u�s��}(��T�o��t~G��S�Y��֬��z�;���Y�!b"4�+c�5]�_�xm�ݙ�~��I��9y�pN�� �.��y�>�qZ�c\���!��6�Zh()�hD���u����G��u�8�c��_��x�:i7�/��6^�e��B�a㐀�{��Kc���"�<�=��s��;jw��{�Y[��
,]�h�n����:����ןo����EAz�Z��@�`w���;GjX�L+�� �B�x����?ns�{k40#�{���oۿ�Zё��q�D,y���-����>~���nh��Ŗ�RӖO~�u%M���8F.��P?X�D���n�E�ye]��e���c�"�ޓP�
:�4�,�=6��\L�/�nׄ�����cS�֮:$��]"�\^�܄I�|e��ϊ3��ܦ2�*��Y!��:J���s1o����������c#�"Z{]���4o�=�|�zZS��La1�N��*�bS�̒�x�t��<��,�^'�����(ų�k�t�I;�(�8U��oE��>-[h��J����a�!+���3>0%3��o�}��M*Wc1��L�5��>b0��YO7J�A4Q*�l���,ō���m�:<�vMh��iCA&������a-! ��x����k ��l���Ɍ�*7��p���Wg7�2N��Ɨ�����V����PT,�)P�� UJ_���1U��|O��p��=z�qD ��H!z�m��i1�HyE��?����3�E��l�x�g�鯌�6o�❢�����@ƞ�Y#�
R��]��Q�&lI�������8�N����9�w�%T�4E&U�0P��Sn��\�C���O�
l�6ޓ���35�Î���������4����1$��!�W��a�>�T��y�u��>���e-;��"���S #���p��Ɇ�O-��S��#��彛=c���Ͽ״����0�I��VE��T���`,���-�e�:ybg-��/�XWn�]�,���nD@DL�"�1����榾 ��c*zO�j���R�!-� ��:������=��sqi��`�n�4����	����`�;�Y�w��"6���
5��y���V��Qw0����H���q9=�SS���G@�O�#���@6��˸�_��[���\6�9���D_�u�=!�P	�ܰ/ns$���s��w��!�2�h���9�Ɵ|@�M�'6���R���E͓��ͽ��Z�.|�����'�MĨGx���R��I������Uj��I���O��l۵�r��q%s�d(�>O�r����0��|���i6k%F��c��*鲙�X�!��Pz2���XE�9�~���Ŀ���k�,��t��l�qe��k���ގT#������4���v����^��+�$���ګ�\��+Y��('VE��jj�Ҵ���rqv�.r��<d%&��9��	��\�ltr�7�������^���vp�`�F�1QP���s�y����b�#�c��2G;¥-�56��φ����d�&�DF2�yx�| �P��ռy�D��{�����[�E��	�9���q����g��N�i�T|�-�3lx�oS�v"����^[�����j������I�S���;o�M����|�\�����J-�2�k��7�>�������O���!OC��3���C�M�^�95FG���Un��[\�W@����H�(��3�J�?��:��+�'>�ck�R����R^�>r ���#;w����*�f@@�Y*�iQ,��t�Pd��`�c'	ԻU&$������u��]��	X�k�kK��E��lħo	;S�K~�	��X���n�`��ʋ�Ƿ���ėk$��w[�ő�DGˊ���T�ỳ=�X�&�} y �t:��s���5?y������$���/ѡ�V�LԨss���E�"]��y�^����~������������GY`�`�_ta���F���K3��h���!")�l�,W�m3g�!�b��XY?Hubf��eky�Oa��r���_0'ٙ�iHZ�F+@2#�֋�(�
���2-`��O�9T6,(� �uʗ�*��b	��k��S�$��a�p�>��}�4Ǔ�:�NG�|�W^+^�_w+0sfA�p�����܍��l9P�	�1���Nz��7�%����X�^̃}�7G�v��#�x��R�>�GbH\4fG��'e��[�����K���疥R\�P[`+�T�����+ۜ��_g�S��b�w]�d�m]�+/3�[�B��* B����y���E|���aei�bx�v��gq��w{�z�3��q�ͯ�kw�n��ۥ<�|п�u����'�bߙ�b�xG����W����6�0ʬ�0X�;�7IWtQ�$֐���	�� �a[�Wa�{��a�|�9�<��૮���%(�����U�#�����o�gQ�����9�8�w����.�O�Zx_�0}k��B(���DZF)��W�\,3�P�������;;W��v�NqM��������£�2bxp�;�P�K{��>��wn��/&M�`��O:����u�(�=���)�ax���y�f�^xC�H$!�-6�0���q�M )���F����^�BM��]� �_��5��q+m�#T�0��z�~����eX>�×�hA
�����gw��ԀHh�q1�#@�G��n�����L��,�". �6؈Na�ORrѱ�A�er���p�����t����  W��8�El�:�A�=[��}:c�6	]>��e���iX�����D8�5�U��/��R)K+L��5D��#�u���{�C���G�-I��gͶ�3?�vc2�i1!�^Xb����~���*�R`6�3�Xd̯�7�, ǝQ\�LX��������gl��M��sUNf�?	%s!�ʎٕD0�cDXۉ ��Q�D��$�,��!�K��,��>̲��mN�$|U�ܣZ����{�s��P�xm�1�xm��cD5�餳�]9�}���u=��hUA��wI����҆羣����N��"�.�${�K��x-X���tϴ�,2I�a��U{��ޏ��yI���8�M�`��M*���m����j����^���A��*�]h ��g���q��r���ΗV�YH��-��?V���t�O�}��\e����8X�e�쉼ɭ�b|M��zm��=�,���Wα���ᢱ�U�tېh�$���Ό�qݢ�����E4�2q��?�Zk>u{A>��pz��kw��-��!$�H�������v� �~p!}�jO�OP2DGp2�+�a����)0���s�Z3�X�^����r�OP�Ni�	�$I� ��|����DLC�݋���<�������� �J}�h�ߖ˟}�5�-M�e;cyAhӦ۷�$8�����I��M/����1yŭ�1�"L�d9�淘��h�BbB�!�D�xYJ�yŧ���v���#��+����N:�m��ضm;�ضm۶�c۶ub��߿���ϻ�f�]�VU�9יs�v'����ˡ��kW�Q���V&�57�;�'�,�Q<��Ϗ�틿c{z[��d7�El�D������#F6Gla!�.gf_�)��#؋@���fBO�P��kA��h����^/2�p�h}.j����W��l��K.Q���-p�|���H�wMǚ��$�;{���W����5��q�(O�6#�/J8�KA�`ܮ7D
v��߿�Vc4n6�Z����_�#�a����[�(�5�!�TǷ,\&s4*�͚�j�����w�D<\��XX��N�j��(8jj��*�����ɦ<�}��歇c��2�`@�r���i:��F�
���l�v���#[�KYX��2��,��}啙��:��@��^���3���]��q�����C�wϥJ�͖��1�Ckɯգ�c{�<��)���~�Gޟ	�Ė�a}���v.�6��#�ŭbN�݊ �j�ז�*�"2<����|UB�E�Z����>B������l��Ly�E���gô�1�7YN�j�Kbpj�"[��.��,�l�� ������(���jj�O�S�e���u^�KY�.U��lb��6�r��nc6l�J�E��|e��Ygޘz�g6���o
��Z�����A9��R(}E}�-��@����zG�J�J�1)�T=r�*�]ln���&u�E���2l�Z���W���Z�b��t3�?�_z�72|�x��K#��6Z�+�@ĕB%�ج.?]RQȇ�?����#�6^sAƀ�>:u����+#�G��\]H�t �W^h�9I@���e{��; fW܎����<���Mpj������J�@g�-�,��&�2?��?�&��s��f���NW|ۑ�'�:c�@~���K�.�lBD���X�H��o�L:ٺV!5�#!�h�k�J˳��tE5.-a#�Vk�x`#A�fO:Dg��Ђ�W���,��hh��U�*!P)��5�]]��ː9��:Zd��ipSczm�����Յ���ӁT��'��a
ɟkc�Yl��k^L�Jm% ���sJ����F�\��_t=��f��ؗt�j	��Fe5?rSo��3��-��a�<�Vit�������'[מ�/�b����aH�6���p�gӕ�!Ӣ9낫L)��5�>�WPp2�ܝ�D[���G�:��Hu��/R��	5�t����]��M1k��RH�zbg%��z��j�2������&�ί�����[C�j  G՘;��ʨ���|N�$�m��ܲ��ư��:��%f �/����S��e�&4�����E��QP�U(�'^�d~��Ϋ??���#�tޱ��]�\��N4�X��H�/.����¾�(���d$���=��~~{����sʘP�����oA����W�z�i�
t6��~���y��1��*~ҫ���/��dv��.d���q��2��n��*%ܛ��Ӭ����Y5����^{?S���9'�fKu1�A��A��Q㮬�yGG���#���C͟�|���5��їoW����D��!*jW��t�i���}.6�w�L{v-�����ｯ��^�����8 ,Dq�Åɧͺ|��J�������d��;�`/��R�D[B\4����(ҩ%	�K���sH?c���Ң��~m�CG��H��*,���V'�\��k�<Rc�7��/�WbҒ�R�tO2��U���w��r��@�:.��H�/�G���6)弃j�D��X��	�P��}j��OaaRh!o(�x9Ҥ��H��A9��`1;�^;Q�6���쮖@X��aύ�3�>S�����������㛝�?%|b�o���<�~>\�1L�����W2�;�=��t5?�%�����g��U���{�f�^��Cv�ˮYH�n��$ݧ�&��0�S4Y�<N��ΘM�P���#jA� �������c�9�;�C��B�����<H�J�p��r{�3��x�\ҽ�G�!@`��T	\3SǗ��X���23��f�����gL�2�1����z{7#?����P��d{^���G����Ku�ϵ|�pw슻_��O�T*�f��p���سys�.��^��RF*��� ߕ�����#�<�P�h[�}�}Ƨ�8a�W���2�����)܍��5��g�w
+ˇƄ�e�U}NИ;<�T��BC�z٩��9�� ���k��.�����9��K������Nͭ���`4��qqa]���"S�+��:���B��έ�u�	ѥ9��+��J���υ���6(��0�^ΉZO���`��_�Ñ��%e�5u���=��B�^V��Z}}�n�jO6x�PY��^�����\�.�@3���i��uG���6��[b1��p�M��i/��JOp�+o�0�޾��~`� �Gvo�O�A*ΟW�#gmNs�d�̮:�,��*t
��'�����F�.E�VH���m9�G>I���˴��	�9ݑs�k����5�����~/�"��b���+&���\$�x�6$z��-�ZRR҇{ Br�B�;{yw��fG*7L��6���e)x�W>Z�曆pQB��M�`4&�}��Xbf��� l.��]�W�Y��n�}���@u!�S{�>3ƽ�ק��͵ڤ�3~q����^6��ED�E���L�k��~8��M�W�Ī���g��IܰRĺ^�уK�2��W*�����_�]�?\5�IN���D�u�.	oZb�z���~��?��P���EUg�#� K~ZP�U��Rl+hX画^w�/I]��By�fEƷ|�3�F4	��;K*YbVG�� �>�R�bh�=��;[h	W!+��v��9��G���Q9';�T�2z6��C��<�5C���zT��K�ܷ���D���-P���e��A9�l���e��J#��Iɡ����2D�����[,�����?îU$����HH6��#�a�������]CHA���|��a��ߵ.������׌��n)̾���{~tc���e�\�f<�����6S�/�d��et��5J��@�}�؜D�k.T<�a.�6�8I��<�q9"���������2��GCM͌�nȮLƭsd>��:���)��C�J�	��Ńڥ�~N��
��qIQ=��R��	�|>��cم�҃���_��c�����ʹ�Kutc�v�	������0xY����@=ד���� a�b�9�F�K,�p$�W	%�QG�;q7i�(Si��� ��s]2 L������x�[�_�5�ح�h3�BA�.�R��T�h��!�$�-;gpڂ�n�1䋠=�z����~=��@��k�ջل_�٪�F��c�!c��r����Wu�fD�}����P���*G@�M�L��ߒ;�D�:_���~���w��yh��_�U����0�9�,)gr�HR$��H�L���7��"d�+%�_pl)Œ�5I|��xr�abF~ 4�э�A ��9�⚨0���÷��f��,y���|�;��L�lt.P����b]Rpgͣa�}�;��ϰef�Q SA�<(�	��K�s��]�ߩ���nh6r��K��:�3V�F%���)ksB�l�6�9�@�EB�! �np�_�[	�$�7 U�s��_�)��͸=:�K��)��_RK���<gjf���a��&�cA�?lЉgx ;9q˅��&�JQ~[�ļZP�����9�}2�����hW�o���?��u�sLM��B�S(��`���[��f�wr�H��`�;�(o�x�����A����na�O��u�KM���5CG��f�*)�u<�N����U�J�~C��t5Q�Z�C��CH6!G�͂�V�Eѐ		}s&	�-��*��QX�����T����g�a�sc?���)�;|*�@�Qv��h�c>����}۱ ��rzB<�l�;��G��������K��i�.g�Iu
���ة��T�?*׷?����SB��Hv�?�'���By�7���V0T8��׶�}&��#n�n.\d�]�����0����n� -w�I(�%[�Z�j$et���&+�^���L��0	�G$�{�+Δ*��NX.-�v�U�ޚ-~k;��c�kmN����'Wu?#,�Us��*Q:�J
�0�"Z�yE�8l|R2���S��bZy%�
���Ke!���pRZђ�S��WB�1,��4�hߕ�VH���(�`Q��a��Џ-�
"���P
�/����Ð[1�� Mdlwʑ��'����د.aE����PG4�,�uĥY��O�9!�/Y����p�
���Z���Ufr%$O��L�RL��"��ߞ8U����}3R�����G�뜨�����$bL�����)��#�_�"t/(�Q���/m�A!�]cPã�f���T�f,*7m�3t��2U��D����I��<􍿇#�E�ד9'��2��#d�+��X��������Na�g�������� �ErPE�O/[:k~DR��4��F(՚߾���{�B���j������O�xopy|V罩��4�索^Y0z�}�wQ/��~����ܫ֢SNJ7ن]n�11j�L�J��ˋ<�K���
o�ê����rK:�j�;�j���iј5/���?	`m
��Ȃuk�2��ۥ�����)�]M-H�i����_���K{L��So����z��������W�)�I�~��Q�z$OVF��n��\=���yvnƽ�-�:W�u.��Y4�y���R�ɲ��x�8��"oB�Fػ�%,�*�E��??-!3��RdK��,�:�6�;K��l/_8]#��Ã�}�.f���Kk8붃-v��|���9�W�KNF>�k�L�<�I�͖E3T˷J%��?�(q�#uh9֡�ى��Lg�|]Ko~B,�1��0ֲ;w�U�bu���G/2+�J���T�m�Y�6E�(�+�@(�U��yi��@I���n��e(��]Q��RL��_�b�hn�7Ew�a*5/}���9���nE�ՓN����V�6�67����G�ݣkN^�.{�Ā�Ҕ�h��9�.�T7����_��y�u;ҍ�b��P��BrD�z�.b����J�狖͆J�>���Y(�����:��^$�]*o��*@�)hwzϪ��{W��q����IQ�vDЈ�*s�	Vb�T�#�?��}2vd/�Ϭ�c�ZM����:�n@=��R��3$F��^���>G[���ס�l��f<ŠK��˪6��6k(��F~��.�`�h@d���2I{�e�LĵXr����:��Y�j�G�-�,�zyz��d��=��]B`&��A��ډ��j���q�K%uT6m����z�+e�m5�id���9(��)�V2�M�aR�*1"����x<�C9	C�/uz2��[�9��D�9F����Po�)}��S���Wο91C�mz�:=�v�ipS��r5��Z�l/�`]>�N12�ةW˟ݮ�}Fu�u9���4^�I���gg��TM�ή��?�Zad�Űa����X-Ew���ydJ�d�(����+��<��g�x�u�X���"V�B��Ki��C�+֞��c��9�l'�wn%+au���|����	 4v���c��Y�:�f�/u:����.�\��N:�'��h�Y�Y=�&�Z\Njrq���׼�V��7���II?2�)�B���M�-�:MD����Vm��S���J��4������/������v(��Z��v�=�<���ʵ�)ҵ�$43n�Q�t}b��##�B4^"F&I(�!��[_�)��:�Sx�!uU�a�u��"�m˼���*k![�dH�`�g!�n�
�+v�4��o�b�7+G�#���*�\8I�/G3����#��
�77Eg7�����Љ8c8�<�17)W+���Ԝ��	;���ߠr!�Hw?��D��.-l)�,"c�%M�`���˰Ռ>H�v����r{��뭁�+�2���>� �i��u���#"R��/ߞN\9k����y(Ҩ�`i��9���6c)��qF �)�a^����9����gBE	)m�
��i�o@$�--��l9r��q���No�t�B�}b�B���G��{�15���+�-�CE��ܹ������4��T�:����ݼ�'���
�.2���VECu9��M#Ak�yC}��}�go����^nU�r
�9��Tv6'ND�'C!f�w|�n&�L����!�&���8a(�h-}`�^�"�eT�n�o�5f�j@"��-�D)�'~pz��`]�T:q�gLň&�]�f�j�9Q�`L�[�@��n�Ɛ�)��aS-�l^E/�����IqyFy��z�	��I�Hq����ex�%��������~�Npr�fǼ� �Ip��&a-ʫ��Hd�����RP���R��(G�4�e�^7`a+,�F̾�&��5�{�R�?{�pَE�����kR50U?��6�0G�r~)����*����G��9iq����_Q�Ub-'2fW�h��]}��]������x�3	�w��e@}W�����ޚ������X�y���Z���$@lL� �R��$�Y[��E.@��
��H��GL��y��_E������tJ2�o�N���uFf�I1|�g�dZ);�Ģl&�̠��V+`H�N�|qx�)X��^=K�U�.��ˌ�����Y�<7����}�1sLOc��;J�
��vO���J��4�O�A#��&�,�ê#lE���E�O��W�X���N�Δ7��Ԉ�.�L����eh'�d�f��k��o�������+����Y:y['��j�9��c���W4o���ڽ��᲍��t�l+ h.��!�,�Շ�߸̛��¦?b�$��$��&�fe+<�z֧�/NH�{�(aB��ˬ�	�!�6)�IE��0�����<ax��^����I�m�쀫J
/15&"Rvj�&�\���674�i�zsi��_+��V��������H%��MA����KK��A�p�0K��p�@Q�Q
F[H_.������XBK3�����ك����d���K��8:���A����L�C��Q�@�**:� Qp2��9��4q	�:�*�d c�0ĀX��4��U�k'2z.%��0��{�ܞ�et�� �4���B������,ʥ��e��ZJڣ�{#V[|�3���?a(hw�tDA����a��er�k�}��$��KrBK��5	o��� �F�۩��<��?όxD�Ϝ	E�\�4+I�9��L+XsBa��l@�?|�
<"��@�h�V i'k�Ü\�q�%��
�j����7��$���H"��%I+�0�5��BY�!h��O�M>$��'����ܚ����.� �~	���h�PL]u������ٯ��X.������O<fX�%=->��bE| ��z�P�6�}=`��K���z �yѭ�;xȠE�t�v���6�����8����o�I1�|��8�ޭ3 ������6f���3��F`�uo�=��ÒfB���O]ݏ~2;`�f-v[2����֊�����)�f�{��S�t�������3�"�(��a��1�b��G��	�g�nX��H�P�X#�Η$���F��Ӗ)*� ��5�ʌ4�����r���Ɓ����~`c$$�0_o���缰A)���a����b7������Д�_Uƙ_:̔�����|� �>S
:�q�{$#���U$��#~AE��}MF��X=~eIz�7rk�`�����z-.o���?\��_#E�Y���څ���;����Iý������� �^)��*y������'W�����q�@�����on��@�-N�se�U߲�+��F/���m����}�NEV��'1��ai��N]��:6�+FN��7�9h� ؝W4Rcd�����J��D\���0�����T�Yy廎_�ߨ��dP;���-�&� �u� �F�����hԪ��i�E#O���'�s�pPZv���\��@ƅC�l�C4��7��Mrk$�)�c��-�
��6)Kt�u:�E�s�~�Se(M�k��X�%��pX�d���\�
�M�|�f V8�"!�����8��/l���)�;���o�����~�]��ghlV9ƝG'���P�L��+�ƭ�,�3�\�8���~3�'�[�Tݠ�N�q�rLp��ֻnLO����m�~19�Ģ��&_n��������-�w�&q*s1����eׁ���`�I
���N��Rc�.-q�����D���p�:����E�l�bڣ�󤴅t�+�!R�/Yf^
�]Z�d����ā���]�e�S�w�K39�H�PsLz'
�X�g��X��� �k�쐷��q�h�Xlݠ����~��J�6���sF�$��&��K����2h��J[�\o�W������kD$�)R}F	�/]�̈́b�B�hA��@���y%\ �aې���TŖ�|ܘ��w���!\�æ��A���Ĉ=��}���׏$��h�|!��T���_�� 	M�1���'d���g��aP���5K^4�����(������B���!ne*���T�Mv���&Zxlƞ�m�,إ���O��As�O��/H��lǿʑd�L� �s<��C%�gl.�o�gg�$��{�ܹH��h/a���I���\1�)�x���i콈�D����Q������6�?|H*d5�]�R���¯�f��w�4�Х�{��"��'o9���E���}@Ү+yL��J��>�r�����_�[8[y�����th>��]�+�^loM��R��}����z|�)m�pE����(��*�,��uS��/'���sfq��S�-��,.����!�U�p�E
1���.�_%1�2_����2p#��p�����k����Z*����E�o%�b�L�Rf�,Wпقcw���\����!�B	�
(�'�` ������6h67\Z
�������*{��2���t�e���u��ܷl��K�\h��ց}�H���	Qñ�Ƅ�l��	5)�њ�[`��U��E�����'���q��
L�J˭�P�O��J�C���)�)�����U \���	*��ep��S���� *L�y���.y�J���K0��Z(����	\�F�=�G�E%@y����qD�vd�����a��Mϔ�ȃl�7X,Kɻ?G�t����r�p���� �g,M�;i��?n����탼�h^��8��9�h�4YY �x��|��"nPPPb6B!k%�*A��,�z�I�E�\+�HO@��&$�<����G}����E	��ֱ�~�� �_ګc��FL���Ӯ��|���y��,ɭ�����%NV6y�@ŋ���K�@N7(�}u�\p�V<��XZ�竰����l��E��9N�A�������gl�gn�p
�'�V��+Ж=)e
�xDe��_ug&iG1{�����Q�
�4���]C���q��Xt�~�� �G�<Rք���M���X�@9��		9��I��w�N�s�D�e4I6łOy	Xp�w����.�W�|fr�?>����/�����W��3�[���l=ͨ�]-嵓U��-�m��m����t�&�.��i�7������GRk>����� ����Բ���bMd��J*�q�V�ʈ��ߌ����O:����k��\��_��q 1���q? �6�g	��R�� ��xQ���Y5>�n6��xnW��x��wר���s�E9���<���I�)<l����ϷB��Gt��0�B\٣��-:�i����o�,4HR5ॱ6C�J\���٧��*nUT��I]T�'���aO��
�/DDL>3�#��N@ٸv�eMq��d�c�����;���VC����ˇ�+���#�u�� uVBh��.�T�����b�h�����>�ж �	���⻮C�6�fǉӔ����3�t��z�v(8��xD�<�pf�{��<,�$�u�Î%���'T݄��sKQ���@��8��l4�)\I��J�.��h�*o<�hkNdZ�X�@��-CXp�-}[DHW��nҀ�L�[�4�`tB5�I�<7�7�)}�J�PKŠ! b���)��L:��h!��ͥ�l��&w�ǨK.�V����+���;8,�~�s�g�"�Q���ۊ����&OBx���^�^_��e� �AC�NЃ�꿤a�"D�-��.��z�c��<aˢM�]��N�fY��?�!�G(Cȏ��p��;�m��'P�[��0���J�f|Ӡ��ƦR�Ǣ$���G?s`0&�4�~dg�ļKي���U+"������$fpH��o�0���`��mN�*�.;��f7}�J?�.s��A���B̟4�E���]v�q����ĐVm[Zu(5�<ic��wnq��yԱ5Bհ��o1�����P�*�@���7 ��V��#)���	�	�����������*-O���ZN��S&��X�ۗ0�U:;����n�,B�]&e�	��1�8'��s%�Lt��.?~���ԞV��夸0��:���J���@�q�Rĥ�B�����."51��N:%&�y���?o�!���xF�k����V�Y���BֈB��S2j����kE������@"�`��� -'��]l�-|���r/I��3���y��j�)�49*�n���1���Ȋe5�-+K��c"L�S+��Q_N�onx�0�6�:=�I	�YIr@[�`2B=��/,v?	&)���s
��n$�I7�;��|#��h"��S#bil�-;���N��S�	���<��}�'K�>p	��O_<	�����ƈ�w�P�a�����r����mЬ���ȋ����g��g��&�*lo�^##�A3�SY��-^�,I(�3�ϛ6�ue8���
@G&�ҥ���k�Ȩ���i�u;:������N��I�������m�L��p���	p���x�2�zh�ܯ��!�sM&��` B#zA�B�xvީ�-��a;���j�h�*@�i�'b���9��^#+�q'+��Ǔ�D��f�z����}}$�"�9�P���-�hSB
s�H���}@�R<&��:�D�ĸ$ں\�N{l2�&��B�u}�a3~R��Mk��B#��	'�?�Ys��[q�B�W�u���F9���I*��R�P9����p���Pv��ݛn��l����0Yd�+l�[��99x�򚝅���w&���ҏ�ͮ]��Um
	]<�����`_�V�*�k��sRǜ�9�}>�y�ᇆ����Ι�W6j�5���.I7�v�����q�×L�);�Sa簯�D�iO��^�PhW��ǥ�Q�u*��}Y���U���#ο�;C��*���yp�swJM�:MeWS躜-q�t;�H}���=t�͊-þ���h:��� ��a,lΪ�)��mwV��5f�����Y\�+q>�0
~G����Y%�M��B�"Ū�$$l���Q�g�X��VC����ߚr�AF�|X���A-{�� �*@L��/��iM���f�E�h�u�����E��d?��7�Q��� �2<��.t��3�i2��?	q5|�PU���tIaM.��@�Eu}|��9l��N0���w:� +*Q�	���V��H�'��%�g,�.y��⣅��}+X7x?���^f���Oo���O?��>���_��ۻѴC���E�#ؑY��i��g�:i��l�XF(BR���Z0d�e�W�.a��=F���q�l�z���A�P��p����������r���Q&|��Qv���R3�b��Zޑ5"���F,�I�chc���Ԕl�z-V�(�؄����������!3�yq�T\8�cMV��U����T��x�2�v}��{rY\ZX�*�S��I�\��Ѵ`���,P~�t�΂V>��1g`j�����^�'���O���y��Ǜ��<�E����BY�K�L|���ǡ\wF�G��u-k��h5.��	qg2���h�����Q��`�s��ڊ׏o�a@���S1���Ÿ���.a��+ t� F��E;]w���������qu_ѦL��|�HK��{�K�]��#�fgU�&���x5#�c���T�@���2��I�����@�ϥ�y���X��Ӽ�n0���T�{�˸�c�xњ�S�O^�O�h}�{؜d�N�週�nV�\��wPd��?�$�8.����|��ޥ���������D�_�8����1���L�f�@ǋ��i��Ճ���`Ej�bꡇ�"]&����>�S�p�k�96D-d����ș��V��L�]�6��"Y#�پ;�:SN@[���������٪��ţJ#\�t���&7q���X��B�@t'�ۺ��3[��<�\���m{������j�ovx���ؘ\_�0�5B�:��^��>U(���U|-�ӭ�"��F����6�W7��l�����4���_��������K�	��-���ūD5sl�FY��ߙ���������],����Ʀ̜:�n���'#��g�J�!8�j}�I�TZ%�#���ɡ�)n������!����t�a��F���LuN��Q«N"�i��>��T#�ny�RO|{:u�%��L�|w�>{�6|��o)���L)4���.���9�z�	P�}�������w��~���Q�ײ_b[�� C���%�d&���'թݻ͈�Р���X�]����c��`�r��9ί�WR�7�j�I���I5v�ח"�b+2�����$F	����é6��epa U�3��	��J��'��bt'<$Ǖ�>�c�*h�5b>6�sVfF�P>/U�_�f&��ܶ��S�����X%���'��Ib�C��݇^�+���6DD�_����tW+��b|��Z�H�[xU���em�`��UدI���|@	�T�&Ye�4F4�
�#mE8�M�i2BrOQ0g�^a��:g^iA����]�M�� Ny�	�\�_�\1T��o�T��z�k1�=���U�&�,̘�H�G~H�<��ߺ�祱Yv?_��Q�����i��=���T�^;��E�|� ��5�Fc�O	$*DU={O���ݷ\�7�ա����n�[D��B�z���x�g�b�1�s���
�B���	���K]q��Ib��1"����(.��zE��7����U�/���o����-,%́�dF���>�i�iR\�CG�+;m�ԛ����{�[�	@V@ 6�1���IT|]���O�K�@�M��	�=[�=�[g�qBbl�>�B0+�'d!������СZ��vxc�����,��5	��������Tb�V�E����OG	]N
� ��:o�U�"ާ?d���S���\?�uݖ#dG�
*�t~���ޓf�"��F5"�p`[���T`���L�J7�Sqw����b����sG�D�|��<+�P�F*����9�nP��D/f.y�rVI��a��!!}Z�y��#i�.5bﾮ>��j��6~sHLB��hk-X�̱���K��Ml�������I�^d��1���w��˥լ\}+M��幪��K����S���p8����p�����bR<xHB@p�\g�U��D�bZ�
��- �bI~�u�V˸���JuPh�-��D��� k5U#�\��~�f'S��d�"2桽,�¹w�;_F��ͷ�-��0��C,�5#�������Pa�H�RVÏ�5�?ן^2���Z�%K`�g���Sg$���c�I�Yb�1b<$��Ɍ	�'���廨߀UR��2��@�@`Fp;��$(��i,��G���x�v��{����!��P�h��9dy������`L�ؑ?��t�ۍ�Y�]~R��
,���7�h�&�%�F]#����4R���c���5>8�yJ�=g�d�D�iPH�\��FuD-���H���N��4x���4���l5��h���a�W{mY`	�R�� ��8|���%!,��+�(\u�k��h���.
Pp�":1c�Ky�wYx,�yjt،�m&v3rR�hӊt�^D@ŉټ��E�Y��'��G�\ �(xKN�.�����8������������iO����`w��5��'<h���wm���AZj���_��3��#���׻\=SX&|��t�e^�#f�5�S�p�0,j!Twu�\�0l�mx����;Z�_�6<���B]A�ʖ4�U���Ebd�Ь�g:`:r����s�|�}����|1��D�G� U'�TSƑ����@2&% ����h&T4f�?���k��hO*�-�"N<8�;d�퓜#�H�Q���xf��]Z��Z�π�#���7)����}�}��X����z� 1B�&��[F�|yf���'j��KV�zK ���Y�I�4%<��8b��PN~Y�p���AMi:�p���(y��4Rm�����h�2�6�Ĩ-D�`5P�<v�I��+�������ScB����%�1fV7�m���22I�ڙq��0�#܆I؄o"M���>��Ѱ,��b��	��7�:��TF���&�K�?�'`��Ϛ�RB<���$��T&����%2���WD��W�cjPg���+(��h��j>�}�i�T��L�p�pi8k\�=g�fǥs|��9��	y���k}%�+~4�L���E&FkN�<Sp��Ⲁkŀ��X�6�[1=k�"��ت-���I�M�4jX�H��Z�F���ly$�Z}s������&��!�C������͒�yS���fA(�	~g0抑wXh�Cơ)C�P�}"�L��Dm�)nŎ�.��] �l�&�m�ZXzЬT�����)�f�j�ns��H�����rl�9oyޔ|N���Cl�n4�9ϲ�d�Xy�T�l\��qTӀ �F�9��n*=��	�7��iV�1�W�'b\h�D��E�p��)CT�=�`�EUbap��z;�6�F0
���@���� U��se�<��PND�`hL� jJ`$�2i#�b�@�3�?�q|�2!�$[������X�"II��\}i�<ʮ�^?����G~m�>�������F����'z3�͂�/B��6L:y��'
�12%@5%y���/�d�%�f�"tZ�4�q�V[��@��KKݴ�t��T��� c�m(�MZM<>��7>���)��r���c�Z�

�+�?J]xG�Tf��YCp��l��x^��цE$�-w��m�q-�I�G�����,�D�M=)��@3��I��^�QS��|�۱�*��,Ӽ�8Eg��]6�G�c�� ��eÒ�ue�_��I���TbO�B��б�i�,CP�x���J��<$ ��,�l�=7{�w��	���`�5��H��W�z�_j��x��.���)JxI$N�Mͯ�hn񲣄�')��J���d��*7�q)���XKC�����d�J^������1��ٯ1�|��n���P���L���6a���4$�\�&�q|Rvg���p� �4W���٨��d��gd�#G�yh�����&��3�w�ї�q�MBWy��(���D���O�'��O�B������1g��f&>Gq{�X,]^;,9�A����G��lj��0�Ɲ�,F��8&WiQ5�ٙ��*����j���	Hh	[u5!�#e�i�U*�^���ů1_oN�exD'�#n�c]�po����J$�.�Q���?���b
��4�]ơI��ɭ����KͲ[0��1l��-��`	;G@�#�;B4�ò<U�����F'�儞�Ql�;�Ѷ4G��&/��u�p�6xG�H�q��r�W���w�?�br��|���1knoˮ�?�@��8���Dr����f|b��Y9e�Q�ӡwӉ�@MV<
1�=/@�!��"x?����?��Ȏ�S�+&�.|�B�Mw�E �d�vS��!�mW�= �{f���î�$o*B{F�\�	~	8Ȳ�Ԅ���F��H'-�,�B�M>�e���߉�"P �tַ`�����tC����іjM�LU�-S�f����E��c�<KiT�yj�g��3�2�F6�:U���s�f�3 ��X&�v�stMN���)�h�>D�X���qɈ��%��O�y��2�Zr|^6˰��$ؓ�Gw4W�m��.�,���d�<*��g'�o������!c7ɮ0Zg����dpE�m�w�,wI������؀I�acmxW��&�H2�P��	H4�gF�y��� �)|��b��ޛ�M��X..���ZR�s�=� e���xJ���'��8 iB��˗�5��A�X����[��b'�F��VM;���u`=��wH$qBBHBB�8~��������G�U���4������-8,��n��K��_�5�k� ��;\������:S}��<U[C]^+)��)��y6����'S՞^g�y��=��g	縓m�����h_�-H֏ �p0�3%3�z��o(ӕ�v�̳��]#N����}z-�@�hi><��r��/����e�R���gΥ�z�~ac��:l~-	�f��{����0`$��=!6�؂nOĉ�B��	��*�Cv�k�u�KARx�f=��Q!�`�/���c!ƞ��q�$^�x���ኈ N�%��/a�﫭:�ϕ|䧢�����JJ�P}x�P�|K0��M?�.è�
M�������,%���u�W�3�����ø=q��A{�_$���$����&�:��q��3eŜ#�� Xm}e��w	�iRQ��Z�� ��@����Rl@	���+�U^>��%.g����p�В�B�υ�0OO����OOV��D���E]�X!�YIG������%���U�	�(����B�=������;Z}���}Ǎ��T�
l4�y�vNM��戺|�L+$��_��:2��~�#8.�񁩾�����b"����|N�-�wX�\�a���f�e��E�52P).��\��M�Tr�O\�`�z���?�+A��#^�~�Րױ��ng�?>a?i�����C��������B���.L����[�����m��ը�V�M9=�!����]��iX�8s��V��>y�}��
�<Sɾ!�y�p�1�IB���|�M��B)��<��a�{���v+#���7�jl'�8������W��������������3�n�g�����zs>���(g���6^P��e:u@��/��M��a��w\���-�.�Y�r����o��$*3�RՒ�'HBB֝X.V+c���k��=�r�Q�dw�Do���ͭ���;E�,��7��Q��ͥP�4`lQ��k�<�^�ɬid�T��ktuW��ʅ(�+Z�.���d��E�Pӛ� nDb�TG�8=:9u��~�)�ڵ�Cg��z%�8����P�zsf~�z����D��9�Րc��&���	OD���ms�WvC��P����������W�]2�s$��Iv���ͤ�e]�@�~�i�P�݄LI)�9Nu��@�h������K�Iq���Kg��^�FV�k8���"b���u�^�3Bո��.��Yح�{��>{EBh�g����P��5���2/e����Ǝ���/�Q����0�R�m��	�ߥR�.RR}�	k�L+EJ��:�������:KC�I�W�m8z3��n���ˆ�[L��pMH�\d�PI�+��d����C+kѷ�9��ݡ�<j��贍��:qWF�d���U�0֒0cR��?;O���^��қ��7��Z��:ێ��{�B)��31Z�m�N:A���˛{��*oa/h�H2Zo"��kH�4�//��j>���Z˙S�]�F0���ղJ�룺<+&����T+�uC/%�7�.���\TbL��`=�5�n�@�ZW,͍����$ 	��;����H�!��<�e��(�[
e��5mg����F��D���v��FI�����0��"��Yi�sF�ҜD�l������^ȾM �l��w,*��>�$p�F���2�����pO��S�x��GL�ק�/X:N��D�����u�h���)Μd���hxd+�t�1�|����iil�L!�dT����aav����THv��	*[���x�Æ�so����f��8�l{��dl99���������������0����{�?��EN��},�>X�Q&�O�ID�Z�aa�P����<�����A+���%ѡ��� ��(}�i��z�y�Qq���[+���&������������V�]U��滵��?���8��F(�� \�L b�=0@�@��7��쫐�E����|��n�2:�)�����cW!�'_ty(��w'B�2Wv�_"[��B��ZF�/��&�-���F`|�L���9�@��#��Q{�0����6'��OLӨ�eYe-{kr��a�V���A��p`Z}�����aOqGD|�s̞�Ƚ0���q�e&;��m���oҲ��|�����|�$:o_�,
�;��Z�"8��r��U�>�0�������8��1ެu>ry�'#��\�j�۞����ú�gg�V�h����Z���J�0Z�XwR���^������7tW��R��2�����Y�=b�K?!� ��zQ'��z���uj����6�r-ǐy�"�(��CV�8�4����Y�3-��^r���Y��ab��J.�S( 4�Rl\\��G�fՏ���%���ʃ{�>[ ����ujzK���w~W�F��=f�J���ΥF��/�I�9�����b�4�UP��J�^`^�=� �u�\�;�볕Rl�g�l_���(�������M��^�f���?�c�<|	4G�s�X�O$�=�۟<M	��y�"��	�Y;��\�h�T�Ud�3�'-e�l��;/
 ��c�Tdk�"�o�;o�f�'JA�����Z��;ę_��p�تD�H��7��:-B?}8TJ�(&QZ8P9B�3��&q;Z�˞7V�v��0����BI�M�.���k'!�r�\N&tk���R����Xv��m������h����>��J��4$��g�����f;�Xy��"^�ޅj�ּ��!��NQ�Xm�Ĝ5���!%&;��cPT�N3ieX;�`�xw?޵ ��yނ�����`���!D�-G�v[�bR��HGf�����T��N�[W8�l�>ѾY3f��0�2����!q�7}�!<��g��AÈZ�"�����2\�Y�����L�PÄ<�]uB�L�!���_O�C=�˱�z�H��7�.k��h%��ާ2���k�OF«����y�ҕ��Ӄ���}@�u�8�V���*�魨Q{%�=�E1�@��M�ڀ̬Ԉ�C���柋-"ۂ�1���=�Y���;�=�8�~}��ܽ�h��;-gy��������[o�g�C��z��>�.�5��� "b�|~*M��i��!�+�<��`
 ���^&��έt�\ꝩ���B���O�wU5�N5���g���-j#��4�����L^���t7˛�7:7kB28�z���ۗ�Z\�3 !�i�cd�:����\l�h�\�4����U����ꀹ��F�W�sW>���}C���b~�J.�W;5*eQ���������{��w`��Wt �g���y]�R��r>^�r�&�t�)݊kO��~�с�����='ov�c�v��絰����k����t��K�P����gr��,�)O��8��,zjG���}��j9VM�S�w̺�������PM�ޕ�m�G��(�_�������?�֑Sf-'���rx����*����x�!G �1|���b/,s��F�K]��͊R��tX=g�*�y��ʂ�����>�%ǝ��
P��XfU���Qs�����y��̑�۔�7�����vJ ���l�&k�+����u3rƔ�>a�����!���Gƶ.-�Tt}9U]"�� {��֌�&r:]�����l�ɔ�[��Ќ5��tDߧk+��_�~�cR�>��;9U��+����a����&b��c@���~��m*��a����q��
`�X�f
�*�E��|�x�I&��j�jG� "��iǬ�@r`��{\%T�n�����Vk�_g�O_a*P0�N�[�[׎q`�[�@�XZ�1�cH��c���ڛ9i�>��PV?C0@���r��}	�I��Bo��*~͘Y�gtt��DS���	l�GwV1�π�?���Afhg$��ܶ;ǩK��K�s��A?f�����|�&��\�fۏ�)����n�R����1�Lx��c�@���Ɛ&ꬷlm�
58-��Wޡ�3t�Z�1:�N�']#:qt�X����ɼrMuSŬ@:�҃��EF�����h�t�]e� ��6���f0��%rY��'�\��!�uxv	��>�JL�:��h� ��9�t��u��B��Ck'����p�:�}����R��y=z�_���`̘���*���@�{NU��$���hoX�;��\'"E��#��~�K��k�h+�٪�����7r+F�~ ���"���4����� �1��h��K��M�cX^y�p�c�<@�@=���Dc����aot�4C $F��1N�L'B��>��؏�z9q��20=��ރ�����r�!�_�_6z�����sm-Р__~����"������u��� ������kG�i~��Fz�[��(A��^4�l>��f�>��f��TH�"H��~���'s5����$2I�*̓���/��fU���<BP�ep�X3��pEy+W6 k��/����KZD�n��9��b�3y����x��5�<���{ ݫ��_�^�ٯ�ٜ�Sۦ;Q
bȰo,�g���j�<@�p��q5>�����$�
$5#�[�+a�s'[�DP��z�b��%��K�k7a(�+��3���x�;�ư��A����`@)��� ��O �h���Q���' _&G1�n��G%�iD�&}�����*�A�*�jJ��ғ���5�����ð���^_'AB�>�X߫���ea)���^�������M�]����O��Tw�RWl*���I���F�a�uةl�.�h�<�&7�9	�
�C�8�q�Ns�	��l�u�u\aǦ�g@u)&?�"5�0����(�Q�� )	ek�@��T���&��J/<.i��,���^v.����-Ύ�o������v�?�xO�K������$c���Raa�y5?ck��ӝ�����ru�	F��Q���Mn���-u^��}OJ��yX�u�B�٦�yJ���y � B:���Y���/� L��t]�"�.��x��p��dھ%�WO���w�;5y�9	 w0w���b�ο��k�+3��Z��\5��z�b�N��K(�4��Q��O_=������d���q�5Pz��a<(3O������j:��t�D�gW8�dRnW��t�`b�rtZ�8���K�3a�u�y���ߣ_i[AX�P8Y@MN��e|���g����T� �䛲�l9jT�~��?����>��q{���}IǞ�J�g	�e�z=h��y������@0Ĕ������̓p1<�]@Ñ��2s� �#O%1�'EkO+��u�Rh��do��eRYl�ԭ׸2�xuo�I��q����W]�a��f/��_P5{�TpVœ��b�j���͖�`�Ig�OU9ݥLi}3�����wG5G�l�.՗츭p)�|i��C�"	ץ��Z~�p!���F����N8�#Ϸ?[2i�)��c���wh��rާ�d�(v�4\Je����J;��0���y�ϳL��%7�Ã��o��55I���k�(?�e�fb.�1W�G�EIHF��"�s����WU����H<s�X��~=�H)��G2n�6Y;_�]"�[2��h�'\��
sSax��ܭ2N.ZOۉ�~���������=>��Ы8�������]�x�H����iʽa�	�G$�jYS��8޾�]k~���d���o��Y�:,�W�$���ֻ��FqѴ���l�ԩ_T�x|�CI��(���7[���\��v��m{��7�P1*ћ%H2�=oSh.�_���#�ߏ�~�'۠6���ܕ�<��t��8j_���Vmu��%�t[��1��T�N��Z�䖝{�֛b:~�H&7F���a��?N-
TE�v&6.��� �x<���0��^�E0�/z#��}p��G�ArK�"s$���7~Ϝ�^JQ�>���֠F Wzʖ���dP��ʺR$h�꿩��%�����L�:���k�e~�&/��WO�گ;�~e�� 48���wQ;�v�#/�^�̨%}�婣�/݁��yI��@�y(m�נW�
f��XTZ'�@:�'�m�xc��C�Qq�#�Ӛ��3L�Ux�o$	��cB�CE���O��F�I�5(Z�����t�%�D�a�z2K���\uO8������(�����>���L�r̝W��3��O����'�e�\�o�z��*\"����DK@�a�)���lJz����N�;"��ǒ44]� 7H��T����l秫6�>chd�Q�s����#Q�{�比pD8�ԕCx(�K�T~��[q/�a}.�y�_��*����FL����F���Ŧ8~���
]���YPbTX�F�0���2rW���w~�B�Kb�rS=�>�~�Gw���ao�N������˘b�`��	�|�����7 �D�0� <?n���d�oR�/>�9ȞH��W.H�O���I3~���y�Y5 ��f��5S��	F�#�c�;���$����4~B�f���BQ"~y� "��\���E��__Ɨz��v��>���y���~E�T��b�S�i?����5M��N��˼Y�"�dۤ����絃�,c�ԣ �b
BHn��akй���df��������T����f+�!~<��G	Fi��7؁���Qͩ���oxX�Q�vJ� �,��� �>4M�a�ɱ~ܷ���py�U;9�St��c{ǩI���L�6�7���&C:��;w�zd􆰧�oQ�.ϝz��,�_��[���Lٙl'h_.���|P�S��65���W�fw_���u�y��]E������!�B��uH�2q�Pȱ��E�%ڮ@�&C���c{�������N��7���Sl�}�K��C�<�Gd}]~	���T#�_zR�%�_}���hl�T�K���}��n�}�"�����a��[����Y��u�WRd,l�D_;a�7�D���\��〭e�?�-[�=���W����l��m��Н�}#gܸ�t��~ib�o��%�F� R3h�}��;w""R"����2D�e¨������E|ҝ�!�!ɣ���F"������M��6٬&������+��E��.@�NåN��Õ6�u��yŢ� ,��&�|C��\�:3���~ZE����wR����7�?�#%�A�䠩mpl~�;�NwQ�m>T]S�_��q���h����������00�f#@�Y�'lGEA@0Rh�+4F��,VF?""�)����ۇ�>�0��ϼ��0q��u.l�w6\6�4��8rI�$%)y�J&ťN<;Z���ϭR�Ŀ��	�N�%� �&s��#��� �+*�G��3*��B��io�9���mX���f$^����g�C�5�6����Z�ٴ�, �Y�MC��H�^L�5'������l-!�C���8F��.�닎��FV�S@�2o���ߢp\��~	E��ўz`/�yV�}!����g?u]� �<_-}^���V�z�!���}?P��g`��W|��{������;I��!���Җ�)�㸊�������q�X*��U
#F�%��a�C�V�=�m�,�39�4��k'|#@���e£��V!^F�,�W�4���C�u+6�Tn"+�Jh����}�ؿ��O�:�l<%u�UÃPtwR����ÿ�T��;��5�iOx'��J��N���x�nB� ��Y��n��JF���vſg:�I�y5F���-�L �"Pw�"2�}?�|�u��e��Hj��Z�"O]h�����'� �&Uh�4o�E�Z^��jK�н���3��Ƿ��n�Mf` ����(�yi��W��td�q��ޘE������[��OA�U7��_�P���T�aY�Y7c�
�2�p�T��sz|����V����N|z���= ����i���c� �fc�&�W�.G@��ut�cwJh��޳��G�ʨ��d�����0��Y�	?u�Ơ��X��'h��5Ŀ~ސMDeAW�̡���hr�|Γ��Z_���lWe��B��MԿ}p��o��PP�	�0E8`�l�A�k��X�dM0�O��zi�������_�]�MҜN�0D�v?)AÜ�g�l��t�IW/t%�܀,���5��c�^rGafyh�e�bWK? �lf������x^�k�e��<w�-��Á&�ְ^[��p���w��\J橆��A�Ɓxy�jb$�f��yWnz���X��j��c�7�s���Lx�BƹC�R�@�R�����t�������W����KQ�G�=��9��$<�7"�<���n?����Y`{Z��v<J5g�ַ�i��Hu�(��I��Lq������=uui���N�b����۸wͩbS*2��N�}Z���#6|� /�U�н�m��)o��$����j��؊�B���Ҭ
�K�R��q�P��=��z&�2y�^��:��0B�<\�Ty:��qs�Ҥ����߮��qr����Ps�����D���`��mFD2��9�d�LLuh���)+~��M�(��A�Me_���n"�W��I6}'��k��TȘ!>Q{i��{!���*�f�?��9��
O�}j�=L�_43�r|iu-�sq|An��Cnυ�rڦS��3"*O�݋:��|��1���*��A_��W��#�`�G�*��Њxl��k�NH��A�����ql6��C�#�Wi�cy��8����N���f(
�Q���DT�ʢ+�4B�y��G�&m9���>�Aóf3����NڠMd\�- -闑��8Sk9:��+v8c�7���%w����I��VT�fg�yUM�e�C:�B<���o�#|Շ]�����ڬ�8�H�
�@!᫖�VSI^�~	)ln�>���?k}�~zc6����\�h�tz�z���?x�a�G�b��?Y;��k��*�2��^Nì���������kc'<��{pO��Q�h+}��of��KQ�����hz�?�u[�ܥ�	�:k���O�3�9&��5���@>k�d�����?;��[J@��|fU����+��CA�+d��f�J����A����SR?ɓ����7� ��̙�C�,Ǫ�[rJ�ʌ�������yK.��Q�Q\��O�$���K���q�O�wg'�����Y\��@^�M�?OQmA���"�B�;����`ny<c-�����%"��3�͝��`:������A�	����������H0���I�3�g��w��!�6�W�C�л�?Sg���-펬۹w���?|�C`���FȺԒ�n����mٶL���2]!&]0�g��O�t$����͡��Ò��������*�(@��u���IJ���Րj(�g��Mss��m[2��7k�ħ!ڙۅ�'�ϱ8�y�U[Y�wRO���Ln���v�q>�۱6l��k���f����m��j��Vm���Rq
�6=!� �5�F0b�cu��V��^4Tk~T���!���\$���?`�U3��e���߇�F)*��R�bB��yjL�(t@������㶮��i��ǜq �,��ſK$'��Qz�M =�&�ft%N���-W��3�X�o�o�u:?k��\A6��Q�B�a@jf*�H%��D��l�?��!f1�<� *rP��}<#r���ϝ�F���˰u~������&kzlFL2��w铣j�tp�cc��[?�< �v�>E�!�D������K���k��m��4E��%�̲��{�>�r���Y	���D��/�^�կ���J�d'���)5�$���I(��E�O�2�T�ɘ5B�`��F����+F�S!���4�o�8HO��ĵ��ѣ<�2��̋����3����5#3��s����7O=��JM�Hy�jү���2�ҥ��g0��Z?t��+ǲ61� g�RH9y��)�x�x�mU��a~:�/1N�qu�`ل�f��O����%���-����{EIH�����+#y+����Y����E�5��3���Jz�b��b6O�{ӟڤs��c�P�&�8Ҭ%�����<I',���؝�𦞄W�M�zԕ��jTc�>&�-B�p��T4X�cP��j6��Y}hZ�L�H������x�0p�E��C�Pe���cT�)������(�5�iUi���d;(��!��	�73�A�����H%��8��eDJ{v�S�	�����q
���:!:�jNQw&��!A���e����"�9ӡ�#������ԪQK\�#hGa=io?,$�Y���Y��.¬"�D��?���������V����.	�E��5����r��H��,������t��FR�o��5��P_rˢ���'#Bw��[P*֥C�`��]��!�G{���ܕH�4
ꑢ�j!�����R��}�s��嵈Q��2c?�;��$��'g�Za��i���_��kBD��}�G&XW�Hީ6���/�2�w�~�ۙ�$.
S���-/�-h�I?�l��+�j��a��`:/��Y��}6`��Q)B�iD!�|],ܒ�D���m�<L�AJ�آ�y�|+KÏ�C�w�2���[.]��4�jΔX��^�6�Ш�K\n�j�7\ޗ>yV*F���&?U�?o#:���[�g5]�0��He�2�xx�]�h��u�&Gf�xL���<�e�L�RÇ��-Df<Ħ��.x�LZR����Ƭ5��ڹRa�ȹlP��f��N_�ъ�dА:x��in�0���*9��Ku�B�l���Q)dE[�>3��MD��|G44�*
�gH��y��Ғ�8����?/.�XCG�yrG�;{�ŅA�=t�$�������|��_F��枔İҡ1��^{��7]�i�&"d�U�1K�l���(�����{����K\)�f�Nڧ���U�k����A�{b6��%ְ�g"�Z~B��	��}k�tbi���uG]w��ĳ�Ws@i ��>^��8��K���]Z��0>���Ǘ}Ј�����������P�J���a��و#a���2]��l!E����b�+�`v�ӻ��SI�|4k�&#o���J���p�ݸ�T�!��k�7ʲ,3�,򇢇31ԗ��!����t�� �����?��L�LC�C��$�Ц�V�t�$T��isGKA��)%�b"?͸�Q���B~�_
�A4>	�u�����!0���tث�zA�ҌCo�J?D���A�6L�u�Q�M^w�r�H)��j��ݢ��`�1�>��� M��
t��h�ۋT��u�36
�1�O�,|�O@K�\>.��E�m���<(����$�Ӵ�
2���"b�K�᷒m���,X���οn[>&���־#��>�bF*�k�\��+����v��J��e$�x�'�R����v��E�n�[����I!`&����Ko[��4Ϣ��O��8�E��C�3���g^hGd�����j�9z)����O�<�Β�n}5k8CZMfѤ�Ȁ��`��̣�SH
���:"���z�����#��RoI')�y�IB�fڙ��3LI��r��L�"K�n�B�����D�W�;C�RVn�Y���S�Q�U�'���[�o�z�ޡ1AO��?���$��B���n�8�,��J)X��5ѣd��wݣ�Jt��V�zJO�����u�|F�P磞��>��}m�p���?78��/z�9�I��N`�H�'����W_�L��.#�\x�����ѭ�Ԏ�T_��o�m���;��Z�ja��TP��x�
�h��B[�	}�*H.��gO��n��9&��E`Ʌ�*���Cʲ�>�C�rM�W��2��O"�����[@!����T�Zf{��.s�,�xz�N)a��Df(?��7^�sF��G����8۩�g��c�<aw�h�e���ݮ`U����2���[��H.��/�&���]��f:�<�7� #����������0իxF�Q�x�:U ב&;S�\LӘz���.L�xWW	����t�dW�?2F��\O%˕�QpV��<�`�6��+��Eq�������
��X7�co�C4�^��J��7nİ�3���2�'�Q��ˣ(�ʙBÃ�|�7A��A�ĝ>�|�LWi����.�<�9+/ *�"\"p�/��s�y-����s�T���x� UX�exS��>l���K$g�^��gH��%i�⥄�<��wA5�	�n����x(>
t��J�4�H?����T(E]�84eR��;��`b_�}��5?��$�?e`����8��HJ�9(�6S5�'KQ`��	�2����F'^�x�G���J�D�'N҉��3z��o=%�d�>3ck\>�wbc�Do�Rs��sQ����[oP���lmXP�u�C%�L�򼘙S?�.�!£�_G��Q?�� �V�x�@N;Y���%a;��H2:�=mHt �z��	�UU2nH�0���D"�w�,�����tX��Z�̀�cثޭ����ߩ+���a99�_�n���g�9+��1�5V��.�p/����| ԒƮ��|j��b�G�{,>*�#p:g�a*x��d!���q�?����B��ΐ�0�Ԋ݇.I�'Y�{$�׆��j�~V���\��l�%B��8T҈�]��~�J-*¼�a��:x`�x��x��b�v	�^��e��x�+q�K���j0J����I��V���@[��o�[�������A��u�v��^�]��<���3�ӪKI�S�]�z��3IǇ�Y� ���>�#B��/9����@�.�Y��v��uK�y\q��?����[��<kpu��`��ۏz�}�eHE��H��bJ֙�m�Y�)Q�I�tב?��E|�bB��.�J�9&�1��	��QӤ^��YCur�@�D�Rq�K��bU�WJ�ϭ��Of.=�EB;�kK�޴	�dD
2���e�~2�ΰ�r_ڡ�0-���p�>\q�iZxO�N�.�Z��AqO|����'�C|��rf����a�J�DG�M�0�TR/lb�=[oBTzt���U5 k�
��p��1� ��Gت!N��ė��=q8�^T�Q�B�OX�vu�z�ߋS��mp�P���U����jJ�$����w�����]>=S?Խ�}�����S�RЂ�ވ@%rV�����t�i���4��hQ�݀3��\%1u%j,����ց {m���jUSL5;���~�jJ/\|,��%��z�j8ܩ&��[�n_��[L_�D�@6PvWC5��rc���#�h����	S�p�$0,�`�e~�5-�Cm�nG`��V�ԈEx���p�������R���(��2�n����7T�p�+���F�[��䔋J���[����o���x�Ҥ�rl\�S���������æCK���Ѻ�k4�F��'�e�ah��A�QԪF�Ư�Y��g,<na��g�f|57B���k�4uL�lz�Ɵ���{�>ۢ��sq�>�c?3�B��?۷��Ǭ3�Q���;N��	ђ��-��+ OK�/��w����11m�ֆf�uu��m�4�<��J־�E��x~�*�j���w�u���#`OX*P��Fs^��NK����{7�*)#�����'��`� ��|U�JA��"u>R&��I֎e��Ѕ:D��9/�D�b:�TZ�R�Ex���a7����E��NsH�}z�R�+X�"5]��=�t��`���ߖV	 �!ǯ���5�0���8By��Lਇ*�~$���&$�Ҏ:z�P��~�����|��\��Ǔ�*�p4Vr2\罹v���g`�􏯎7:($��p{2�k��|/!o|��>Wۃ���5}Op�|�//P��0�tɃ�6�\(��W�ݙ�f1�()����xZ�4gT���Ћ[Ur��S�<���� �_��Rq�RԔRTPzʍ:mC��I���v)yt�h���r��N3�[�šn
�7�bS��UPx��R����<�ƙ�>�~[4҂��\	���I8�_z�T�z'|o+�[����)L�=�Y���Lꄽֈ�<4�Q23:&�=�r}]�}ؼ�@m ���x�t�d���g�>�J$����ŭY��C�R*�N�g����T�#}��ҍ�?�"^[
5R�y9\�����������E���(���A[�vj��i��[���h�nv$��[�x+�������7�Yʞ�bW�EK]�g��梽0\�`5�!����!�'�b�������,�y��gĭ�KgMwۿՏn׈>��8'�z��~��4�|�Ц�_�_��u��(M��ЫUې]ʆ��w�9N�m�p���d^xN��8v-�G�oχ�m����9��^*�֋�/)#2g�ئs�a�AU?i�-\�N��L��$��š�c]�\�n��b6~;�!�r���F�����eCZ��^�
���6fA4z�2�w����ٰ��P.L���(��?�D�{c�o�C�����(����x
���Zt��P�ה󨮺��Q*���x�����X,�TlӃ0���Ëw�%
��V��Ǳ ��g#`���'g7���#����$C�;qwtceտ%.y���o��5��h�}%�6ɭ���~&�'���j��V&\{$�)&�S8-�M���U�G��O51#��Sp�~�?����ߢ�fڴ>.�6&?A:�x$
{Z�"�0�RX�5��q3%��Xθ��Wt���W��`��s3Ka��d��
F��J�0}�5������+G���� ���!w6���cݣ���l�4L-j�n��vF�Lu	����Q��N'���-�}c6�[d�Y*����.��p���əp��a����8m׽ӧ���1�a�d����d�7�夷-����Ѱu3?�����ɢ��%���L?U�^�#�D���F�aR�[=�y��d����EbL��L?f�<�k�!g.�����I��0'��������xT�a�/�_������ϻ/�E�]k��]�3p7��3�JS}��7���C�-��.+��9�$�mX��.���7A��)�F�?|�	G��v��-���/SD{-Ŋ��d����#���.��D�����`�@3���6|���P�y��闀k�Ӑ��:�䓱f���]���g�@7>q��a~�f�m*F ¬���~*�j�ڠ���q�^#��C"�m���*���w�ڀ,<񀷰h/D�ʗ}�N�3i&�P��C�V��A�L=W1���9��pȆs��}k����u��y���g���׸��*�6/P�m�>��<�#]����5��M����=�L�F%�_S��%�֚xM|���ȅhe�R�$F��G�Ô~zXX9�|u�b���#D��-�w��/���u�QgْՇ&���w�)���Aو�ӊ��a������X��������?'�»	�r�=�
�$2�D�s�s��P�������P��)�g��-1�A�j�v(��+Q�;.Q��"l]�
���� ���5�ޣ�aF)����@�]	���&:��Q�K#1�����!@���(i!��>ߞ��n�K�Fum�Y����[j�u,aӈ���9$T��S鄮��]~x����B�C4&���.Xu�o�p'E�� �_u�yG4��]�%UZ�Oѵ�u/���(�ε�ꏉ�@�]��
dL����δ�kO%C�m�~K�z���/���Tv���-�2|�cvk�p�t,%٦�-�0�oԥv�:��ӎS����*�AY���k\��8aJ`�ZA�2�t�2(
��4L��p�ͤP�Qd���~c2=I�G�	E�P�1� ��F���Q��{�9���D��`F6Mj�@*��/Vr��7׽�b^�jH�ȪP'�@(U�a���4�>��^�]��#�N����gi=��/��͟�+�-�KU��V�~�4�zcӎ6��\�S�$����7�Y����bu��I������J���:�g���f���D�&8�.� ���=�����J�	�q֜`!|7P��{+=�(���-������r�S%�3l/��Y��2�o�@ts�ӡ�p�^�*���`7��૑��5Jl�(d=���$�0�'����	�@B��r?9WX噎���;+��&���V��p�� 9�T�R>,oP~O���Q=w���(�_�QYBAY+�8�-Ӱ=!�R?��I"�{���(��t��ߕt�]ޡX�C�#z�,����<K��<N�M&w	7�؃���O���B���9�	χ��Rw�"g93�g���s'|IN�F�Ű�� ���}KM�"���N�������߅����_t+.���p.,͝4��t�)ƍ>��q�$�����fn�{�.{�]!z�\�>-�UP�t�r?�Y�$殸f��ޡ�g\3�C&�m`�yV��H+NS<�v#�LRC�M�Rτo93�d�/�;��E�d����7���#B�{Q�c@�%�<��!ƺ<�ڳ�}�C��y;�(� ��6X�?�?&�9:��6�ضm۶m�۶m;;�ضmk��%�ﭷ�_}�꾧���U��n����,���qH�L�[�D�3���k�H��!.�Ȓ�� �onـQ����%eoj��߉9�d�:�qi㚤g�G=��+�c�T���c�a�+u��n����[W��~j�Ҥ��/�ܦZz���n5�i9���j�L��r���2�u(�Fr]�/�W$l�������(O��<�}Aq����D�����=b]�nPE��qit汅F�����X����l�z��N|g��٬�Ž=5)?h�~���۪���?��|�Ҙ���$F�]������F�t{"�C!�o�*D�~�>H3�y-� ;r����~,1GӅoC�b��:+��ߪhF��IG�1��20y�,/B�T�qQ��ZEK�it��ޒܼ�[�H����������������	��1y���''�M(�����S��,��F�e�����A����ůȔcT|Q��Ԍ�
we$�q�1��f��� i�=���~�C��=��8�U�6�UR �`�l�o�`��gN:gR)�q&�f�3�t�y�����\t���Zf�=.�|�'��� �дB��t֬�+�P�(��᚛9~���'�����h����{�����k%<��Z����e�k�cv>fGfTs���V(�ꕢM�n�@�P�*�y��w�3��i��C��;��u>�<d��羞�$nw#�tw��@\��Kow���m��U�`��ރHJ�k`T=a>����65]��O��c�+y0� G�0FR�����ޥ����S�Ɏ>�������j����9xΗ?�k	(��o��7���c�u�o7�g0)*^�T�X���篓Q]�ڡ�����(	��2�����"��T��@];�Y�*ូF2\����-��.�2 '˂�J�}m��R�����VĶ���D�'*��~/0��;��=�VpĎ�/�BY�������}���k�sl�6�B�h����Zn�KSLA:�N@1Xn��-=�zJ��Wjza���]̗�k��D��ـ�!���[��CH����7��Q8#75�K��a_n�-T�:sf8K,ٻ���V�O\�@3�,���ﾴ�Y8zv�Q���M9T���p�B�B��D�&�;��\�oޛ���/I6����d�}�݈d�i� Z%7�6�8���=pviϗ��Ui�OV�{>�͝Jo��k"�؟��/Oݗ�#c�;kY9gKy##�����L���" ,���+��SGr��ۥ!��"d&�!��핀��q��#B�ގ`���.�����~��]&B},oy,6v��>���5/W��#CG��H1D��jՔ��ws�dG��2�I'%IU�l�K��$��XO�oV˔!&j$��.����:�� <M"8S�"�1n��C� ��ʘIqL���z1�\o���ky�a�8��k;Ux�.t��Ҡy�4q�.�I�+1+_�b���=��ڨ4@�h���&#�B%^����w]�=������M�y��6E��tm<��abEo��D��3$�0�h��N�B�d?��sܘ�M�����r�'�L�c�Di��JI�sQ��|bI^ឦk[�4�!v��	{����)��Q:�feg�j�X�v�D���Hqv$�M��ޫ�v8θ����`���Ŷ�A�Yԃe���e�n�E߈�r���Pft�
�#d�yj% g6���Z2(LQ9��`�����Y�q�/�9�-���1@��&��9��;�5%��~�Dπ2���?is)�� ��q����]�pZ�v�w~'0�H��Z%�q�����)��xH��I5���Ƕ�2m��V�zZܹ(h�U�ڥ��8VX@$�Ѽ룦���b!�1:+5m���;v�H6?��k>9�BC��	}�p�al��I���h-I7���:��N>Ҟ0�j�\Ӊt���g�Ѐa4�$����|��]:Q��Nadc����.�)�nj-��M�W���@��L�0�[NZ����0�q9AIЏ�n����I������rՊCH=�����X�}��b!�mş�0�AM�U�������1+��ɥZ��ʼc�&�hR(hІ*C��"�iG����
p��t�,8ʄ��3�P���_�K�-��"��~��W�������SN��g���N�s�gfyY����m��Q=�����[E
e&�q
c��q���������E��|���j��+�A���������N8OiV4� q�8�T.ռ��C?\7�9����nq�[��@����b�W,j�'��eɨ���[s�š�'ѓ3s�0*^o�Cܾ�ѿ3V�Q��'M��X���t�+�(�:��gy�K�>kAu��4)��Z��J=E���t��������%�O@<Lq@�'�#������'đ3B�XC6\T��e^m�,��� 'Jm��*�N�5�Y�b
R��_Ƚ�F퐦5eTL�RN�0��dku��<%��;�m�#�.1�P����4cT����Fqz� #�6*Y�*��P�kq�`�dTC~���.#,�(C"�8���ך�K�����ݓq�'t�{Pw�_��7ǝ���b6!�G��J ��8U�R>�*�YG�1xFQ�ZYY�Z��S�E�U2�˘	/AL�=n4���#p��H��.̛�Ƶ�=~­ͨl;�e�%�-(
Y���[�X��c y:5$f�B�dbN��(7�u9R�����p�5攷�"N�

 �*{Z��qվa�1��*&mu7����Ph�݀[�`��{:�����,�����B��Y��Ԗ���xu�z��ܼ��!��^ ��T��(�('��gM� O��S��a���il�x.T�r����Y�����Di�g��e5�|�
�d�f�Q9`1�5*B F6ڏ6!���X�4��ǳ���h|2D5r�-0u��[��]����G���`�=�](%\�רު���$N
�����*��G�4K��K>��Q�1MW(b��""O�#��HR�u,� �Z}�~{���|_�¨S��"��u,:��*�r\��S�����ĺ\~�e��|�f�˖�<��	���e�R��m_� "�EC� L9��!m`�*�Ǧ���f)�]�	�[!����V����}]�s;?D�'L�H���Eɺ`'ߓ�/�+s6(����sLC�&���\���7�EW�A%(���_]���]t/jN����kty�9���������G�F����u1��xuDڷ ��W�A8�<���'q�-�Β�V=�L�q*�`T�10`��g"1�c?��r����Ո�\�Pk%�v��dh� �	�V���-%BG�t���N��������($� ��z�қ���o������0J��S{ߢ�����c���~����a�V'�I�׹9ܝ�ð�����_�Q�g�rɝ�+&e����|�F�)`�~{�V�1"+|:��gu|�m����r��v+�u���.G�,$`�F�k��A�jE3�{�,8h�C��XX91��9?�����B������s�G�^Xem��J#�r��n]��ψ[r7�WD�{����@��sr�ڲM2<��t�v ~�&،c4g�D��2hl�Dn��Λ)�I,C<UC�,�����PĔ{�[������ ��宷�y�<9is6��5�j���!#z.�M<V*��������C�s�F+H��XD�I�H���#L�a��<25,��6��ṫ�>��ϊ5S��X�ȵHk���o1�ySO��6h�%��s���D��T(���.{n�v�i���{�����o1�Mt���A��KN����xM������``�N��gW�dا���Aϖ�h�ϗN�����)'RZ>:8��I%�d�`�Hm7���xI�x	��@��1ǆ(�c�� �PI9凣�d������Rh��#�m��M�_����7��x��Ls�*�𑃊κ𯮣��9�Q;w�	�����tF�O�|��W&��5δ�>�H�.�rBHL�/��#.��,�rH�*�j��~��k=�~[��3����b�sn��$� ����q��p��%�E���=��S0��[&���?��S��K�C���!�+��x���ղ\����
#��B�]����(	rC����gN{�R&�*/Sf�=����(�oG��-F�VC���-���7ש��6�"���z�~v�� ���g���Wv�����:}K�e��M4��������R�:�������(���Hi���GR�]Ѿ�ES���o�F���5-�̟Yoq�j�ɿJ�ԕ���/��&7ת��;����� ���B��|��ܞ�����z��^����e��^<g���� ڴ�����U9$h�@��G���ӏr�ODEy�3-��O{��[����I����rۥ#�U����+��-���+ؿ�/EP�vG�<�`&�#QD����d��Hf���4*�	r�h$�`�ic	C :V���iz�K{���nk8޿���.+�c<�=M� �?`�2"��{���h�穵�����Vk��G��?��ė�C�¼�M��!�ܸAJ���ZˍF����3"_��#�+$��KG��cfx�+R䝏&�}�vX�cj�S��4u��~�.�O�������!u���S{/��-7�����S������F�̜����	PsG{���P��K��2m*?�_�<p#N�'D c��&u-�;26	R>ye�>4P��3G��S%iX�txz��7����&��.CX���6��5��
F*��>�r;lvev�3Cm��@���@A�X�x���[!}�-����+��S;�IP�S�,��^�vv39�o�pR��3��ٲ��DX�VYT�⋯tB�������\9f?�>#YЫ2HXӚƬ�J�[86����Q�>��A�k[g���l�,槂��(��}��\���=L(��Zڇ�z��~>�^���v���`��p��Y���	�@���)����S�Ad�{�\�Xf�
mj;�||�����&W�{�g}Sa�V[�6��*�r��ըz�֩JbQ�I: �X�1�v��s��{9�����K؋�	f<�C�:&�z�tz�6Dl�2d��b��,`X�ܧދ�~��у)Y^��t%���6It��2? ��lP߶��ʛ��	���_��~"7hh]S���(��ww�]�{a@�� ����C��a�)aŰ�j��;12f �V��t_�d���s���CK�����U&d2��y^�w��îȜ���ˌqQ�p!�)��U�%�#���G֬|��&cbzy�@�1v[��d��,�!�������4��Z.ױ����%�H~ �Ԭ3�Xc�^�N�D�=��_ë'�P�֪�4߫�� h��I>��a�#�N"Ƽh�t�����'}��UÆ�s���̕g��]�5�i�*O���0��>0��F�#�`��\����/6�)2(|��{u�_�8����}���~ m���#����BG��x�6�~����K?���q�-h�4�g��WY�f\���蠗K�r���K�vt�)���SR6c��ӛ\E�z�q]'�ŒJ|N<�3w�}kƼ�'7#r���Z�s��3�S�b�S׎��c�k5���,�
����m��^L=\���K�(Bi�q��&n/{ˣ/��)����#Nȕ3���^6 ��^2-��.�ר�h$i���~��D�~�:��'���a@y�u_�C1�%�`#�ɸ"��#/MjN��`(�I����9Ҋv�(X�)����o��銃��i��#`|��ĺ������D ��m�*�bR�:����>�s㥑7b�\�CJP���9�u�%�^��Ѵ�G�kԡ��jD���}��g�. �\w�I[�Ҕ���vS��`&����4�~R��W!���r���DI���f�z�� $
�ǘ���P���ϵ�?��s���b����I��-֙�Yv��9�
g��H��Ŏj�sA(5'�'�Ux�P{�-�V�j/�ʚ�ƙB@gi�<���}`n*K� im����S�4x�!�n"��wۣs�5ܣ�ܞ��M��<�G�[���)n��9:F:2��k�h�\��ɶ?��-�Ƅ�сL����|�2N+Ѡ��KI�����:���㭪���co۲�me����@]Z�0DYOX5���
���NNʰ�$�IX��8."qPVn;E�OCQ��H��p�u�)L�1�NicvU�����7+�5�9��Q<�#FM%$ƖJ5�3�vy�Ԭ�ؗйPy��?\�3���X�<E6�k��|)�ى��}ݕ��YA��p觴��R	�j�����9����C�;F�i��
l�<x�:�l<_ˣd��mO6��N|�����F��w�Ƶ��'�/u�(���Ո�ۮ^�[��@G���o$�I��<�RX���z<>ʤ��X�}P�uC;��t��d!��V3���e��Vj�y��̮yw�8�?����#������ny�gg�{��I�1O^�d�u�xx��<�<��2��5Z���� ���D7�� &&�r�S������������G<I|�z��)5�l-6so�+e��4T0[��ġ�ewo���0���*_���Ӥ- �u O��8���Xr�ꏘ^���Z�f_�z������V0�P�tz6o�P���0�2r�sˁ\LR@9FY���Y~�p�h�Tw�E���h�#�I�D��rd
�#zpz��UY��E ���Ю#稖�6g9"?�cQ#���a�F��l������6�N�i!������I��6�HD���+,5/��s1��`�5�@��X%�3OaZ�a�9�S�[T��(�4O[{AOr�3�U�v��q�N�#%"j�\1qFRH�����l_�ֺ�iUə<�{��3=!~/%�=�zl��ꪋ��A��������o����_�����E�ш��B���O~��N录�ե2�u�PA�Hc�)Y�'�da_c+ً�Di�]RsG����b���n�G��fV�#�m}�	��t>$a/v�69�X��#4��#�SRC!�,��_5�6=n���Z��"a,�a(my7�y���㲵ۼj%@ķ���9L)�����_�����L^��I��2�úe`|��%WΔ���tǞ�P&,�p�h!%aү���nq�K�Y�w����E~�M�q�H�,�\Fl�/���U\d��a�����ƘҐ����+fb��t��Z�'^� d�> b��p�tg���69�,L�_oA�O�0���,��,,�w���Н��A�fᶹ��:�-9����N�� Δwp��m�Y�>�dIr��)�|JE���Ysh����s ��b1UKʔ��D�9B8���wKry����O�
s�0�]����*H)qLa�w(R�n��6� -�f̼�H�,��W���v�a�m�Ћ=��tJ��=�1�5r��m���� "�2����Rz�H�g���ZJR�h���`�J���)���"QS� ���ׁ(�l�E��H��_o��[w���4�b(	�'�����i6�;:*�TAX+���Ȉ�&�ɟ���\=��U��x`\�x.ȊS��BсR�sT�f���������WtT��N9*�v��+�j�}v;Bq�nIA_���v:9~K�����@�F�Z1ĳ�
��AjH���|�NT�t	���w^Ů��Ns�rh��JT�ܧ<hczn\���K��A�_g�G��KT� �[>ET |���YV�%�&�A��hx�in�e�͎�@}�F��[Mo����o�.ޝ#h�t $/���;�F���w"��n- O$K�^Zk��_���Ӣ�C��k�@-O�ӌm��K��P�-�k�+)�.��_��B��`�+���it�E�P���pP�{��L���Z��E�Զ���8�
��Ц���Ǔ�T�؍�A��owoW�T���R��(��N�l|;;0j/�8��d�Yw]��#����u���]
��$�~3V��ڥ�|\j8h!��F�G�/=�����M/( �x��/&�k 5=^�79W��"	:�B��<<uR�C�C���&��#$�'��b�vo�J�����m�B���߸�ё$E��)R|

h�k�GE���8��z�8��#�*��$��e^3v�|ӽ����m_/�^GK%>����J��$����E�vW������TG� Ģ��IP��O�A�]f�M�s�ûrN��w�1�Y��J����a��t��]�ݨuM]\�DF�x>�!>�g+�%����ʬP��ʋd�{�����.��Ft���W%�0�,�i���2&�E��Ƒ�6�VL�O ��|AWL�Q��8FH��� 9��\�B����ouMP\<��>��r���kfbe�M�
�[��%�MK�UU���^/������!��r�D�k�M�N��{n*�El�B�
bgD�V3DT��LJ�dt8l�-�6ۗ�c����].ԅ+��e�����]�l;�<�)gͳ�Z$�7g��]�7�j����g� 5�&��
�����zj2c�MX���osŒ���0�H1����`�C��f�Cn�%GC�蟑N����aX�F� ]�J�e�c��Ki� �WgQ����]i@�S�$�A�9�  ��b$N�������ֈJ�0/f�����UϺ50�i�r6��ީq����iV�=��'�	��]��]��;-z���������a_�n[O�o�I�{Q��Wۤ�9o����\Rufc�˦��e�෼]�ؑܐ��$�F�f�x�r��'�=�M�s��9_�6(z�܄��v��;7��넜g8l)��%jc���6��c27�կ41H�-���%�_Z3���=4���4���+K�~����c/����@W��^��x&L�)�a[J.p�b�fZ�-�C�?�9�*Ž�Ff���f�{���Hnż?�T{���Jo�����1���v�����Er<Α��<"Oh{G��Ub|8J�Ʋ�5#~�I���ࠤF`K8�g3`��w1�-
!��˶HMhmҒ]�D>(�`�p�q�K���������_�O/���Y�o׺��Q�,V<���CY�:�CB��B~ڜB��'`�幤���._�8�a3�	����j3_�0�&�r�u�ph�o#/ؤ՗fX�%����7�y5��S�`�W� (�3�YE��J�l0H�K�f��{ pDn�T�q���_U����-�:3+F���慽�p8�5.o Qr��9䏰*�/F��| �i9�A�J\l�f��x�MU�7Q#Ƅ�K�P}���cmA�^6��X!=5�~�#l&�\M
p���}�B�lJ�{L�/��H�Ƶc;SUf�,ޤM�ê�dW�r�2D7���ۓ��C���Y��{{�x?g@�0��в�!�� ���ۃ��l���Y�d� �ं~� �@���"0걸s��ɨ��ٽ�Wh�$�8��G�L�)�I+�2�_���w���i���ѿ���� �=�W�0CeR~!H�lFT�쩱'��Zt+i	��D(-5�*��K�~�16l/���N�Ha+�$�𚽳4�"a�<,���2j���P�Y��j�!1�0��d�q��4��kЅ��{��3'�Z��4�����,<�`��G��bU ���О*l棑>I�f�s/�]��ʤ�A)�W�0c�L'X�eЪ�US=<�ɾ+�G�ar=`O~���X���H�X3!U_�$����2RF\d?z�$����L�O�@³��d6�=u������C]]���o�������լ~$�.��"�����UF��&��\�=��p��U�n����{���Ex$l�P��7$4��p�n�_:M��T��R\���۬M�3FT�n�}��)����O�:����<��x�R}�[YS�o����ǟN�%����,�$;��e�� %�&[-��k��`%�K�wg��1�l<�,��Z�
��x�Ur�
YHEr������#Ւ�ڢ����Ł�J~���p���x� ,L�R�������~K�xH����!7��(�7"������`P�� ��ls�������X�9R��k��T,�U�a��-�X~!�%��Ѷp�4�~�=�.�����2���ARb�QS�ryq��\�2l\�3��Թ�B3k.���t��iB'�MJ��#��{�Oc C���(7�a����~Hp� �8���q�W��gi��Rۜ�Hڰ��Kƀ�Zt%����oU�4�\]:����H&u;�g�w��f��������Æ~ğ�k�R�0�,���_RU^A�#J��~g��5�$������-N^�/w��E��_� �T�?$M�YrYī�@��#���]��,l�Ce�~��- �f"��DA	",?:�@4o%����"]۰3��b���B���f���P@�/6��9-y���ц@�C���Fe�����D%&$��"ٖ�-^^���.�X06�i�(g{�>upNy���;%He(~Ch�������G\�����S0���,v�LnNw�vbN�k�C{�8�l�Q$M��G��M˦��z�>�
���o:y$=!>��6c�y��t`=T����x���7����TZ[��ےZ���R�!P~�%S�E4��*r:b��?�-w�w�h���挠��Xr�L�Ɉy?p�:��&D�(�4��;m����kW��	�a�
��@B�5r	��NK=�g�-����w]%j^1�0�W;r�u�.X����#���˔���?�:�x�g=����Y�v�3}֞�0����N�ܸ��N������,�6�c�a<(b �BYbB�7{�q��~�7����MdP7nB[n^�Z��in#j�E"���A ����>l߽�u�s��0��A��l7����M���C/e��}��m���VP?c�V���se޾Oz}d�~�m��s���W�w�a��È������`�Ȭ0o������3���IQ���0F�"� 9/����p�+0��{��H��V�A�&��\��?K4�p�]�;ٽ����'�u�/�!�mD�7�D�W����y�߾R���w�X�~?�{���b@e���������}���j�wR}j�U�边��e�l����07k"����C����Wwf�F ��9�1��g��g�da�qa8�5[���e��iF6�;cM���n$u���^�VI;˜�,�*f�~1����M4���qN���bdi=�꒿~*<�V����\��˩�Q$o�X�X)
�BѾoż�P:��?"�2���`���0����G$~X8��e4pZ\U��9Xl�}U����G,�Ͱ���%�'��7����ťh�$!<�&�2�Nx�b��q7���2g*FB�
���8�e.ܙ���������^�^�(f�`�SW���v~΅��T�9���΋]6~���4f��}(Xլ��o���<�3t3դ��h�;����&O�ⴍ�.�����z,��T�8�8 �<
(C�g��'NK(B����M�OtAb�@H@�'x�ϱ�170J� ������Ju�6P����н,�Cq�����G���cZ���E����u�7��b�J��x8�T������c��%�&l�l��2��1��Hə����v#Zx���&Ҧ�W!�P��(����;9�Kˠa"	��ՌD9@#��h��ҳGZ@��.!��'�H�5Y��n�3+3��A���6԰���e@kjR��A�S���w���
�8�2ª�ϸ��<'���[�o�Z$�ŽMB�?f�@�t�W�i$�7��s��9�x?�3
ʙ�+�]�m��=��ͅGUvi��67�)bz�%nG^�@Bπ��^Ɵ� �h\�Dz�c-��v���D�

�ɥ!l���/��vÜ7%[�6���G����k��/f�ǂ��k��*��悲�~m�ر�g�3��*���H��+j�t{�)��v�Xgxf����=Z���,�
��H`ξ[���nv3D�e���1��B�\=v�����V
˖�?��H-q���,fg�	�ф]lٯ.Q�E�+�� @,t޽M�,��xH���Փ��|�`�b�g �an��z�|H�S0�3�/g�nW�4R�!�ͺ�ɢe+��@�덪B���{�6gټ6ohj�kf{ߥa^��/��C�r'(�$t&#���(K*���qk�y3��t(�_t^j6m�8�uj������h��2	C\%��A�"��� eŐ(w�����K̅�ˢg
g����6���N�4��>�����y	��V!���.c��^AJ�_��q?��
��Vzϋdo"7�w��+s�/��캛~��ӑ猆�77��^Ϋ�iN�o�ߕp�eZ'��S�:���u0pċ(A�s�Q��b�k���fD�����T�(42��eT"2�����ұ�;ۊ����RNp�y`��D/��Ɂ�kP��,� �J�i	���r���g���a�r�5i7�h��Kk��iK��^���i6���K�nx��f��Z�@�̣ɵ��i�f����R�Ķ_n麗�Mn��U/�x��������ە������
S�b�8�I�٨��O5�Gp�pF-^f`���)����ezP�S@���EW_��9�q����n�u@+�2�p �����`(���|7Dw@<
�`�b���z;�M�h�6�Te�z�v�4]-�����5�
dN�=g���<C2)i6yҲ�$�7�m�,
A�d�%�0�e�9=��qs�0@FS�O8z�쮍��#�]�A\�MX>��%7����?�:}n�Ɋ��б#�T7p��vv�
!�l{�����F��ȣ]>�3���J�E�-��^)�&7Œ���J�w�4���$�g��!9y�@�f��e��o��M8�d�	�s�1'�j��$"7�M�l�Ē��M�-{"S��MO ������T
z;���j���J"���z>,�`_�q��%Ǥ��I(�R���{�֖(\Ǆw���M�����Ͳe\���H$ �����u�l0\�)����[�5���hUP,^��Cеm"�Rp%�*?�d��<m�U��\��؝�]�C~ZH��8E
�UsEYqy �5���Ib8�]nh��i�مð��vE�K�(��`�����z��y��?}��i�51"������j^4s䔔����gU��V���7�zB\����� %&%;�,Z��
�IQ�QR�^���̲x>)���cx/kZ�^�߄�u��=�����~kBi���[��XH76\oi����Z���s�Τ�P
^�<ct��+�R�
���F6���4I )�C�,���v��arcI���[��/�n`3O�=�hs�O���
�[O��/Z���a9�Z��1S;I��s�^���r��fY�$9k^��	��D�]��F}gy��01׬�_����4��?X�JmBU<�+r�>�IR�S���K�p��덣X��gn���i��5��8�XO?]{ܸsjܭJ�zZ�8*�g���s��Q���wjX
���JZA�,dC֔��ˆ�NPQ�Dl�J ���]xpR!=���.?m�@��,��L��]����B���-L��1��q�O ��G%W�P�^w��֟?Z��ïS�L��
T�����e�l�/�V�*I	��ϬXE4v���Ꝁ�U
�A��ڔJW?�#�UT-JR�(S�`k8����y�YvhE�Q��J���⡷��+�������\V׆�_+�"K �R�ݜ�5?�T>Z��Κi?}z���k���+��;��'���;�3�C��t,���0"Vg��W��2ϭ���u�u�����SRQ��d�u�#E�|����GΛG�	ܟwÄz�밑���xm�{�ޭ���������(.�Z���ئ&J�'��0_;Ĩn�Qy���X�]�,�Y/�*�>��xǧ�LD��L�@�v�^�&4���K^��%b!�:�|��f=3��7�_c#��$t�����d�4�.B!)���J����	��i.�/'As��q�)�V����Rw���tG�E �_?5?�f5g�?��n��!�?��^���VOw�W�T[cW�!E���z}��x��J��z�LS���T�s o�$j��!�ܤ1zE,��q�0?����4���k�<��25zy���޸��ۂ����h�!u���T�/BCpD׆f��_��-�bE�fO�<��ͥ�
�p�bd�F!�����T̹���E(~�h��Vx�R�k��޺l��D��C�6��5�	'���Ͳ67ͥ���s�L�M5W���-H1��qo�m������Uo�I�u9e������9��AN�:���&^�Kk{���G�����.Q�dk��ls���7�Nk�9s��dx��N����)��xpޘ��s(�� �����e+��ۚ����h���u3�ܕ��_|��J8*�/��<���=94�ݽT^r�������sy��"ʲg�H���Q|o"IJwV��K�k˪$g=�B�?-4�ɦtx�C�;�om�>���[����uQ&�W<Tuӗ}/x�P��,�G���˺/�*����7������}w����Y��bGrW���ˬo�Z����e�}�_=���r�_�_��'8���+��
%+�����lev���=?��=}�r�Q��QHc�,G���iħ��i*+JҖ�t��Br4���䋴{�\�a��~6��5hyӻ�O��B�.LB�� ����s�3 ���uIS�����*�a�B��W�1�Jk�98��ns�|o5�<}S��*����ͩ$���ߵo����EF���[�fsX�&�"�9򔗜��ⶀ��Z��C�=�/�ۣ�4����Xk�߫�<���DT��)�S8��I��i]7.������>)̥�F�
�fJ� �����/(�N��ߙ�@�S�7|8�׀�F�k��t�Gbj�ԧ^g��MAw�\��aԦ��d�;��Jz�̡�?�nv�M_ ƞcE�@�P��n�E���R.���m�S(�ʦ��/���~�����ER�;7H66�o9e��E'����(��k�M�@	���:+���Tvyt���n��N�o��e6��s6p"��	�������g貼M[B?�+\�a)����9G[��e�0�A.�y��-�q2	�W���x�2P<ݭd�m���ɨLv<3٫;O���E�&ɹǕ��>Їܬ)���鍣8>��L#y�U��ǉA��܄�*�,J����� ꉱ�w���?�vw�=u��)b�;ܽ:^.h�dUN�/��g��~?pY ���b��s3k�e޹��8;9�%���|�h�e�AG��]ݮ7���)�ڡ�Q�l�����扴~���wF��K��Փ:ImA<���w	��&��{`_^~�!�d��DB���g>J���Hqx}��h�5m�i����:�Ξd=�J.����	CX�^n��(=�&|Dx>�V�oYY��ߔo4�f��S禁�3�R�1��k��f��܄���U���dr��0��zb�a�o�R'�4A�����Tc��.t���^$�d����s�Y����r#���]*M4�b��E; N����0P:�短����y�4EƆux�bF�f��@��6���rW`M��g�%|��N{����Ō��#p)r�o"-P-�d�~{M!���᷆�����u���[Qd������sD���ԸwE��#�?���HZz��e�����#h� D�i��������%:�8ߟ�n��dD
)w�+.8=^',�UY]�M/�D� �X	�߬qt�H����ld���˻UX33=��v��oó�~`��
������ʊ�����ﺳE�QT�G\����"�ﺏے��멧a���'���(��O)2a��ѥ�&����u��oG	���	/8z��H�f/^D8rJ�,�CtO6qݎ=��8pj?�e�]8��~d^�Mh���c�T&ٛ�Yz��NZ�h�Z��Ԑ���`��{� ����Z庥K���a������e��x'�t�f�:��w�ůH�_�Tn����E���.��$1�������8uӕ��7�����\6�����!�Ns��=�7t�Z���jR����QҮ_0㋄�8̲���c+��ʋ_�5�9��� *H領��?eF@����8=�PT�z��s�O�QC�D�`UKu�obJ)Q�W�p���0	����]A���Si��u�oy�X���[�.q�&�+e?�E;����a�zBI2��T%Qh6z�F���do�ƃ�@!����V���W���M��*�>/���=-���s���i�ủmN�m�Ll۶m{b�۶m;9������������t?���F�ӛ�>�M^j+��H�dX�*��D����P+$$*��ힳP�٧l@aӭ�%M�yBh?�,w���H�Ԣ�:h��|�Omr(��-s��Cԩa	b|�8�����e��y�D���������0�V��|[1y���Lާ���Ck����I!�f�[�ع`#׽B�KL�UB,�H��y��(�C����Z��p3v�ͅ�bIr��_������Gjp��>@����G��f�Q ��	�m��%�6����?H�v3�����ϷV�M|w`�Nmx�iL�d�!~H�s�8?0¯��ĥ�O-?ǲ1���{����*ݱ���Ert6x}�p/[��V���X���[m�jX�w#jӚ������N�{MZ�:���
��mϥ�G��~r^.��/E{մ����Wɋ��RI�鍄x,�2��갾��W��'��-���z7
>��Xqb&ߗ�R ��٣�F�5-�p������AꭖV�]-� G
N(7&Կ�H�|�`�L��q}�ػS�^�����s��6^܏����Ktj�g�ئ]�eF��f�J<��R?v}ߢ|ӟ��M���"��#�N�����+���[����y:�_1y�lÇ�
�vu4Xa�>�|�s�?#���>��&��n�e�F�b3��2�'4�\. �����?X]�mw4��N�'�\$��w��I�_�تZ��aL=���2>��kp���L���,��8r�ݒ�Gz{3Ӷ����(I%�?�E�����!��=uPv�����B�'�Hyyŷ���>W�����y�>N��ۿ\o��#{��]W�c�i��J����?i�ŝ���T���BR'�i��O��}�0��.vʝ`�^��	#޶�d�q-�5�tC����#��*)�{�|Zw����Y�z#@O�qlfz�)�Lk��S�;����lp��Z܎�zzJ��U��Ud��=�M�O:���i�#u,WB��T���d��nf����+���M����#�B1J�aJ��@xO��<���N:�]]��^v���a|ۋA[���̠�T�z��͙d�m�L RcR,,4��f}�vSB�ݽ�Y���t�IQ����z��fF��ґ���i���mi/�p�L©X�JlD�ʤ,�&����ҥ�x�|j��� ��T
>־�@ �8�R#\b�Y�{n����@�����Ec��Pn�Xx%lA&�l�����"���0�/�-��#��|i?۲��#mtغ���#nxM_�m���깮�6��-�a@zH0jcK��#��d���K߽z#�d��������!x"����k�K)�{WI��љ��`��3��k��}z>������=KP��^R�̶Y=ݒ�����#�အ�y�f���|�b�Q"�����c���$Z�|�C��)y�ߌ\�-m�-��'S��4A��R��E L�,pRC�a����b:��m/F���M*������xͽ�78�7f�([)�<Ne .�1_@�B��T`PX�U!+c%��@�	F��quD�`)��Mg��3Ӏ��JϚ5^�뎽�p/�J�Wg8��J��֎#/~�<C�@T�x�e\���A��3w�c�t�;\}���6%�8��ۨw�q󝶸���_�'������,5Z¯xD�q��Hw;Yk��|�vHf�sb��e���rj�����$��|�W4$��W/�(&�?�����>���h��{<w��E7�5vO;y%�/�£���&� W1<���
�R��_}�N��l�@�!d�Ҡ�ꗆE�:-Ur�9c�	Sy�F�٤�&*I·����jIƴ���W4�>��CJ���N�2�T[�˝UYz,`����9cy� @��r��l-��G+����ڪ�s�/�Ő Y �G1,Z9�㣜P��F��p�?�ĸ�mfH�Wj����z��i�5�t�5�)[p���OO���E�D�W��$�x��̢�!T'W{�8��d��aq��oG���U��2��Q�1���9 fy��va�k�����o�� ,YR ;Ǒ�%N�s�Myᒡ�`�-:7��}^��Ш�՘��0��2�!��m�=�7�[`��^<̟j�5�S�N����O����0��|50
L���B�8!����R��}��F��j"��穌�[?t'�Ϫ#���?�Y�q_8TlCם{B͗=��V{y
�7D�������9�r�b��ؔ�M�(ɉ������EVq<��< {�l`��~�m'@�Qp��Z0Ҕ�᪝�:kK�̀�}4J��6��j���@�Ӓ[)؄w��f�E�{��n�� �,E}��Omc(G^E�P�X��A�ݵ�HF��JV"r�e��Y[vS'<�uA3��p#y3�Y�>TN���$�X��n|����>E1p�JWN��?�CG�B���=+^n*0�I[�/)�Y���5��W><sxNI�����~�?�TUE�NyQ*ϰ�̵Fa�\���A���)�C>?wV��YZ����ސ�EX�j��<�RC��Lx��1����zzY�4xz��~�pj^{z2,a�lp��e3A�y�೰g*���BO���4��F��,x�4�91y��^��d=>�5W�XZ'����׭l��g	@Mh���V�:F(�?ј/�O�X�ײ���}ø����ל��8|��:�+ٗJ_��ӻƌ���3yx�	��㸴pɱU�<��������S���o�p"�����{.�+B�/<�m�R��_�'8~k
�U��He-�T(�W2�ɗ��^��(�z�ہ��f�\U4%�jMe������\+��Hx�]=�"�i٫+o��v�Nbq�6Z!��uV)?Y�UΜ�2����!� f"vl ~��TFn��r���V`�W䧏�h1>���4T>�K_����;�2�ddC��lFՆWx�S�f!�f��b{�wW���ko��5�Ad�����W�'>j69 Ku�H:)lIi����G#4A�&��#�3�'�kkX}S�W�"$O�|ni4�NDvD��K���QFPP)�|N/	S�HĒ{�t��A����J䵱�����p^k���ۻi��� ��a�O�_����$m�;���n���:��(mG�6�ܺxԩ�G�;�g-�FƁ����,�m��􏩋�ǈ�0o"�<�Äț��q��p	���8N�B7Ȋ;��*�!-�+�bj��L|3B��؟��ĉQ�B�p�5�*�//�F�J
�Nmow'��9�盝R�?.�(:�&$z;k�����-L�;zA��Q��v��M�b��-y?t���
y�j�}�CWg�Ǆ��?��#�p�K�y�sU�Tr�W�K��	�>H�펝:PkyU��+k�awgf�˖$L@��©t�=���7JŁ��B����l?����B0����@�NN�
��iW�'r%y1ҏt���?hT%�� �7�R�ԑ=��id��-���������'�C��#����y�=|�5ڲ�4�R��!V�bY�es�_�eP5ʑ�22r�P۽�ꉹ8A�x���m�͆%_!5�T0��}�.��un��^��cM≎�#�2/d�Ihր�rf2Ir��B�A���i�}b?�7�;���>���|�<�q��|���PM��87榥�q�mȻܨFTA3�q:����,�A2�����lHS={���p����d�8er�����A�Mv�=K«L��J��h/��I�>n��">��f�T��y8����,�Ĕ@�eJcb ���fti��*iٯ����K�@�3�v!����xy��S�OOO����>%�����IU�ep�'[>X��̱�0�[�iqk��y�� "� �2���I��1��\1���]�Jw�Y�e��M�FM�	xX0�v��@�E�9���<~��%9�L�<%���D~^8~J���a>�����Ԛ�*#c��Q{E���rD�VJW҂_N�"G��TEmgW�E9�)<@@<�F]CC)�M�
9����қ�MI�V�ms5����<lB�Oy�0ab�(�x �{Ϙ�ӧ.)P�fo�W�OP��0��,�����T��+΅�w����4T,�*o6��~�m��,�/��aS��ex>0>W}ܶZ�Ź�f}P��~s�vK�]dY�j�&���hzJ� 8gT�ο�+�m�uP�N`�l��.O�p��4�CT��!d��;6	�:�hZͬ���G��rTar'tC�,��u�T*�j-U���>x�ˠ�
t�K��}�LWQQ�/oW�+�:���OӢQS�^q�B�A��骣J+����GgF� &(]4J��|i��`^�lw�ν��g>�����9��Ҭ��Q����%+A_�*|��4��B�<z�L;���n*~]!ds���ӡ�][��Y�O �*�0\� ��?R|��+(�M����pNҮ'��ۉ���K�!J�5P�e�X���bJkI�p�T5UiB#"P�9��pl}���=+ɘ��;�J��(�ڤ��\!-�kAb'�1̩cH,�,��$����t���@�1�nT��*jו'�_MW�ryTQ�mn�u3=e��.M���k፡��tǽ6�DQ�=��㯝��"V����lx��Rqi��T5���ޤ���h����T,ށl�����JQ��;��;Jf�7�1η��D��z�v��k�?u�.`31�N���?U�q�f�έ<0"�nI���2$�l ��	s[�3SfԫT�{te?���,���$p�6��&sM�����4v���:]P�I(��!��ϓ��N\�|_Ӧ�B�Ӯǅ,�'c�����	Ms� �
�S�(���/#���6�i���J#wb��ŵ�w0�onM�BTv�~u��a;xъS+XFr��J�r�\M-u�&Gȴ�݊��͞�c���~l@p.A�hwb���q�6�u����j�9vEߍ?�i���c��;�V��N����qd�pN��a^����=_! �rE����T�2�oL���d���N;¾'^2�����S��gcb�Y!&a�W��zr�N��+�D�$L��>-�&�=�oq���J�:��������?�!UN���^oI� C���KB�N�ga��ب$Fa�����y$)���9���A�^Zw1���A�
R�UT��r�*p�8A##��VD�b��B�FS�X��)A���P=�dg��!�ʽq���\�)�}ce4v{�Ȩ�:*O��gH8Y�4*)d��d���Ec;_�KGb�Y',YE�67��[l�R�Rk��k��|}_�~���W��suńE��_������W2Mf�'V۶��EO�,b��vС���)59u���d��	Z���>�u{QS�I�5�g�CfF���q����~f� ��f�][����\i��D��9I���g�q-�{0��*t��J
ѯ���?ɦ���>pX<J!�A���z&�Î��$&���G��$Ėa��(B./iP�B��f[���
y��6+C]Ñ|譲��5���g����\�^��G��q���%�����#QF|\d
~�絕ҋ�Ԃ � �"��<�����GX�I{i����@����s�m+���3�*n�B�Fu��H,At�C���H�e���T�,� #(hux��LR�H/�G;|n}�3�֙�}���E�ƍ��(+WB�ہ�!m��<L�Z�.EKKK]0�g�G8e�/~�@��~'��l8&(����%�q7S@bh�zRӎpa�����=��2��
o����*跤	W�*�.^b�h��G�/�!3�g*�8�1Wu|�������S�0��ҍ�+�wJy9A����K�<���rP�2-w��i<	�a��Z�v!jƣ�3�P�}�P��>��W��}?�锚mA��pY�pO��5Z�"�@}4..N��\	�X�y]�ow%�g��.��d��Zג�TP���g6�<n�b��X�C�d��F]ni��Z{�i�K�G#cZ�-����P��\��ϟ�U�\�K���{�롷aU�X/��s�|��T���
Wɗ.��z�@�_3�שF��0��
��b���6r?a�M/8ˈ6��
}x�1 �V����"9�����^Ǉ�ф�$��޴MI���S���W4�dH��dO��{#��ԱG�6��9�N��?.QJ׻X#U����n���ˬ�
bu&���C��4o
Q(�\��h�|���n8�j !�0�f�����c�宕ϋM�4Jo�r�G��j�/�Y��̟i�p;Uɩ�:�d��]ܙU�ǧ��]LBJ5�x�"���_*�u�����f
?67�r����d�!�t)�'�'�-'T<>&q ���
�,�ɕ�/h:���W@��҅0�@�A��k[��˜�lEiP"7��4k�T*���x�3���:Y�Q�!W���c���$����(Fu��eyRtQ�@�ۏ	N���~��|+@��y��g|�� ��E�jg�E��^�xrj�6	F�J.�jA8�-K�Rם ��\���hSմ9T��eK�(bD���V�y��,W�|aMd<�˶s������XP��eT/�Bz�A` `9���Q�p�y�t���ʖ1���pOW�Z�c���k2s�?8m��Cr� l	��ș�`�`Ϟ��.S�����Y#�5�Ţ~��ҽ� P�T򉀗H`?xw�/��arI����?�[�ʡ6���|�h݄�7���)�)��(�F��='��fJ�|��JP�+0�8=�j�������Ƞk�b֌�^D�*�"bw��loΎ"��i�֠`П���q�� �2��g>4"a�È�2䴃�wG5�z�|�����z��N��[>�Ȟ�b�	��*��%􋬉���{��	'�N�U���Fٻ`dْ��)5r�nL�#X��� w f�xS �%��y��6.3�!����<�����h{��\-(��Ϲ|'&.������Y�l�<�Ka�q"����Q;�����t���Y�A��vbW���BxK��~"����!���ɚA��h'��֕}_iV��^�q���l��#@"�R$�q�wZ�pD$����f�8�Tep%`6� ��yA^�"�"v4h��������S^>��h>5���	��J�jS�'���#[6>�0���?�V�~�E�geGd͔hGY�vڦ�deVl��1Zx�vǙ�����z�,�K��$51�Y���v��=�HƵ**�󄫺�|F�:�=_/ή'�@E�*��D���j��vY(�ꚕ���(��Q�,uM*-�Q/=p������zZ�t.�C��|�*�dǾ��*_t�"��֪nAa5�-ŧՅa�筱hd�)�5����ŠP�	�3�M���ew��ˡu��$�Ax��/�?A��~nq�6�و ��0�>U|��#o�왮�y暏���H���V���Y��� �3i���Ж�tY��cG�]F����(��F�X�ߴ��45ZiB��7�&��Ⱦ�Q`5p�S��`%ͥ��ֺ����>K0Pk�{3M�.��(T�71!N��}���\+�5�;��Xc���,�ْw��(�7��k "�p�Ⱥ��{_
�y��� ���7 f`,�m��1��=�}cS���u9�e��A͎J�$8��D�Ư�;����~6�(����
t2@�1=���pb���G����ѱޜR����a��L2�S����h��i%=��y	�nac8�:�`q�Z�B�Yѿ�+9R1	ޢb��|$�)_��痣��Y6o$&�3���J|��L�7�i@2.�v֭���c߁�06&����{�I��O�Q��}�@��Nn`��_�|��h6�*��!2�{`�S1ٗ�@����wd��p4���Wo� J�6�쉌r���\Rr��2���~'yH���B�`ӎP ���%��j{۝1�� 	/!�����(7�%�>�4��~'�ӓ������9��)kU���\g������U���ht��K��h��ޏ���:��qۼ��I,�3����g	;b��FS�A1��kJ�W3�GW���$�9A�1*I�!�TH�-�ђb��a�+#�54�I$���91_N�i�jۈ�U[�Bx%�ֈ׶�������R洕��4G؉�T���t��L�2��SH�* 0M�TW�:^���/�������/���I(F9.�<���"��\|A��<!�"�R?2J�gӫ��'8q��)��I�O�1K�^���R����c�O��c�vd���{e���ih�⾛�?Uқס�p����%�7���*N��,8�z%W��]��m��\-/㲴\V��Y��ˊ_�D�r��赮�%<@��E:�NTt@�&R�5P{L�a�ֵ���ˮ%�veU�&��j {�s����O��v.ƃi�%-Bp��M+�[�R ��ς7Y�J��g���ʃQ6�rX�,]%y\�-�O�i-����7[���=]�Rd(�c�{w���?:�+��g�Z!�rE���G�!�	�hU�$��2�{%=bY��x�~���@�t�ޚ^ij���r�͋�s5��*Dp���[��=�%��b�x	��AS8`^����5��M�1ɟ�U�����:��#��'m�u"ov��RP/o?���GO'9��bl-�� 2p�^��0�W#	}L��8���#jq��^H��Hδ{�a����{e�����P���-$���I�?1o�/�0��֐��j�ކ���������IGgj�Yqƴt�I�F�ޫ)�%�o1��K}���n)��v>�v����;��\|��]�07�|r�D����or���Tv�c
;�a\��mo��.����gn��S֚fd��pc�?4�iú�S�P�Ȓ]�O.��|��Ye�F�o�UM�{
5)���>�E�*r+e#p��?���V� �"`���������>Z�zἫ�b��-Ee)�3��օ� t������X�
�frI�E�5|���-��$Q�����4ljuH�M8"_����t��B�Q�4F�٣"�Q��:�5|Jǜ�{|봌���"c2�{�&���S�F��頴
9�uY�Js��[����>:�Q0/�ZY��;
�N�&�x:yI��ʤ��� V���i[�F�¢D�cm ��F���krFf������q��L_+eW
��E I���igsci�����G�Ά��F)_��?+'��7'��T�Lr���!w�5[
f+[�M�/�A�@;J���6 ���j���+�3Ā��*yj�$�DUeyW z�6���L��	�~��ށ����%
O׷�m �t%X�(�����c�%�~g��r�	q�Fh�/��z��O�t�QR�,��z��j��:�>[]�f�`����!RA�Q��j#eyZuP��t�>-�K�/�+td���-�ͣ�Fe<-�-��A�,rD�FXf��Jܗ�]缛C����������4ܗTF�H� z, �ʀP��ul��TzQ=�����k��B��a�x��J����BZ|���Zz��/3م�9��,]�u�<�3�%���x����˞I��\f�e~B_�.�\��q�2��x�Vm�h���{�o`��&]��O{wd|�k���E榝*��	���:8�mG���%.P�3b��d�E�@YT�	���{*�%���=�7û���z���%��0c���?7.�����Ciu���5�i�N�I���e�d��5<3#zW���ŧ�PDq���I����j�-P�3+�4�����~��9��eֻu�oL�����tt�5��_u
�쟈���)��7�n��u���1���@r\������ŋ]�������|��~��|1ё�h�D�:-Y����E�/���ݶ��t� ��ܘ�z���������G�6�#씍�p�Ѡj�@Y��3����������n������D�ύ(�~'lJd7�nT�w�����}�H9����Jx���H��܊�v�b�MMFM�ߒ��r���-���F��3��^2�
��������!�PT�ʹ}�0�����_(^b�"�$���!��1�{1l�N��L�=nq#I=ʰ�������y�uvꂈƫD�^�u;�F��|=�oG��y�]�6===�@�x�z��G9@��^T�&� &,�7Rmji�x�g����j��������X��Q�zJ7�ȸ3к��/`���좬��ߋq:������nq��z�n[5>d!S�/:��ȱ�� ���n!X�Ť�.�՘T���ϔ�I�Z��#�2�8/ܑ�@��f7�_t�O��YW����ʝ��R���s���5��7����Ȼ#+��?���zMn>�
5���{0S����uj^#��:���#nIy���&���0�����l!i�[89�{q�g��Fߦ����=�N�?M��m�h�G���Ls��6jp�ٔ�|�Y[��%X��6���5'��T�>��"0�G��"|�e���6d�wѿź��/ C��n�?��&t�����@����F͝���A��J� ߯�i7���	:N�/��N蔹��KN�z4Y�!���j(|��<I�"n<c��x(�׵�z��=�q�~�P��G�(5�t���G=�S�,G�u
�m!�3�/�x'ZH3�BQ
�^<?"�0
|w����U�F[�8����Pu�围\~�Ɇ�f�id�j	���i4^�%vϥ.'��3�J�3o�g0b��:V�N��:<���4������/Ψ��C)�39ϋ����p�-���$��)x[��KF��Xw����r~ m7{�`ڽM�G\��p]��)|c����y���*fi�^cӫD�l��Ȏ_�B��J*�K��w�m/P�|+C�\pK:�/��B�l@��t�3��4~�)%!c^]����T��4��&�0�c@g�����GR� ��W�]�b���q��+�H8,)�%���N53��A�8�lU3��F	��=�"� CU�k����BP�`0����;Qv�G��*��a*+��E�F�(��W�s�̠cӏr�3�y�[��/@r�t�;�ۈ�;tn�SR
��eJLN�+)�fM�snãK�՛9�7d�6e&������E!�� �4�Q
q�wN��S�[(Օ���7�DV����O�,*�6A�RX|��J�wr.��0�����f�d6xѨ��*.'玜�a#R�=��M�e�!Ii��ȫJ� �F.5%%����� R�Sk)!,�Z�L�=4�B�Wʩ1���|]SQ!�>==�3uzO\}D�̐>�t��̅p�<�k��ֽ��p#���}SM��o�u_hZ�j=6������G��u�!c�X�x�@l�� 8VV�ݵ��6����1n|v��̇�&��ӯY�qƎcn�&�>7Wy_x^��� ��gd��era8�����2���#\�
R'k��B���"���Q8�V���V A	�H��?K�9��#��8Y��51xI�CM�c�mD謷�����ۿ����v��s]t+�m�g�X��_���?���<��%,y�����!l���&#%%dd��ĺq^:wf�Ə��
��&"e�ۛn�h�얤��*����V.G\e�������E�_��/<a�i��Fmbe̵��ab:��B���8�����b��0�����N����k��.�B4V��F|��؞���(��k��ֱ� �z�z�TF��U�z�V&��=Ø8�� �e;���&.�TZ���_�i���5o�f4�����?`&���j ����Ʋxp\6�L.o�2t�j�����Q��Q�K��66�n#�9C���"�C^ �э�`���|��t����t�˗׷m�;�>�'����7�C��ŏ�F��������/'eK�z�LLL�%AZ::��喔\�0��j�

E�ň4�64&FL^������!((��e��.� 3�\����3�/~N�@��t�>(8ѷ8�� ��9ϢP���:�� ǅtN��/�p2��S70�fl��듥,��A��+��z(AW(_��ڥ����pO��d�Ӹ�w@}=s\�@�RCC�O�y���=�\9r{�xh�Un�å�!W���h����8C$kl���o�d�]nA�[��%�^�]=g�2�bCUFU�)G��+�wG�-���EC#'�L�o�(�X�Q�A��e�?V��S�!Q��%�o+��}4_�ʦ��E��aq��D�/�
�R�Y|�=�{<�\t}zs��P��A|��iu`����ϙ��F�Xh��^]f��6�ݺ�����f!�z!��Z��a0x�W��;�,̸(F�D��M[u�)A�k(CkI	���9͐�f���l%��9
�s�+�ϭ�M�JP&-�I�a���`�J����^
�66�p����.�����n�w�GA8.ʰ���<���d�����  �I������T��HE���>v��=��D)j2�0Ei�8�?�	)$`ے��I����B����ٯͯ��<�25/淺7��`=3UE����4�qR�EOic�Qg~ǡ-@�e��K��x*�.v ���h��r�/��k=���#�Q(�?bK���!E����Ѣ��O������܋���+W�Wv�"��ӹ��/�V�۱_K�n��iT	���f��@�G8rw�c�n����>�b>����{"�ɰΚ�k���-���HH��a-���Gʜ=J5d�a���>�Y��,n��52y�o13|<3;��[βX����A��4%�E&��K���<V(��rScT�#���Z+��=7O!�Ŝ�Z��0�{��&iA�*���M�V�?S�: T{�y�&�/�({>kchM��^RцAH����	Ă�]�BcA(�ŝ㏽�Mм�<r�$��&����w��~�K�ș`�$ڵ�џ/��#��,+ۮ�/�W߬,;'3�ǡ_�8�3W##'�z���p=]6�D�ւ�nj�sI��u\<+�B��� ��7���a�py�9����E�ɻp �����d��}Z����}�muv�/&��S�>�&���nك�iYvq:h���ZuR����H����_��pX:(�^W_{�bweww����s���ɸ�$�`��ܜFX�Q���]Wa�p�
Qsw��^��_L&�Rj���M9yoť�	P-Թ� �>�z�h��
�QQ����T��ٛmA�^�:qO3:q�N��T�m�(�K����H��Ǒ gj������e���4E��-��ǎ�7�s!��䔔��]hdٽ"$��Z|�#����.��`=�{"g0Tu�B[�"Tz�\�R&*x��5��e��W-Ggfjoچ�f��y�@���?8�d�seAi2h�4�{=��k�{���"�p��t0�5��c� s^���u����f�Neҧ��.�_6�"<������5�c��i�7j���2��3> w�?�<ZU]=����g@A����#ӏ޻��f��|iZ�:�[R`Ĕb��J��Ϋ���U#�e�8��,ԕ��zmə�UOO�9cz}Ұ�Q��PR[Rv'����c�C���j�wx�c��ޖA�	��q������&17���+�h&fO�f�Tgk����E��z��c۞c|�M��b`m���K��RK������0�,~p������W!#��+�)�����7G�`"tI�'�agI�
j"]� i:�V��t�6 5v�3�t��ѣ�>O|x���5q�mp>�GO�"�6Ջ�����"�|^
���_޾L��)�+�`��#,?��~�'�PlJ��g�=8�b����/S��a&���)��E��:�����g烌��-��n� ����Mǟz�ERK�^\�4j�=�mO�q"PA	r��>��>��_.U<8�?^��q�����Ç��Tp�@��Ԩyi�?�_�>��K��:X�v�2��Qg�𥞻J| �`���o�z��s܍�w�Z�F��h��L�g�@���lTv9M;�_��F�Y�i`q{�j���;c�ȕ-�y����p�Иa;�̦���p��y=o�{�_�K��/X�V�3�N(�����`�����ah^�dɢέһ�ן�j��3�E8�;t�+1Lf�_|�No��$��y*��E�$�[��fP��o_���}��aza}{:t��p�7wUR���=sv"A	^ɪ'�F+O�JV��Q�%�<��W��h=L�)��i147���2�6�v?0/�@Y	=��_�R�^�ސ��OrH=��Κ�`��md"T��t�W�@G� tbY��l�R|&���5��k��a�:-}�����"�B�v�Ek�n�a�{%�l�X�ݹq�6��FɾAU��HOS�W���i��|�׭I[�� -�U_�(G��2�q��?�;��7�ƍ����������TSK�!�̲A&q�Y�M���C��ZTJM����	]�V�]5��m�ގck치��~��,d��*�H����Ç>a@����T�§��g�3�ȥ��	��'1?Yz+�|����a42��'n��?��VE~�Na�f�+���;{��z|��@-�$NtV����/G��o�ⱞ���o� �Of�د�5J3t���hF;�]�_�<�233o�f��$Q=A͑�~5xhY�N08l�}I*���zsק����c�;��Q�ϳ&�E��H>�!8������.��I�Ux��9�:�h��[2�?�� 06���1� ����0�ɻK�1��-(��<>+E^���P�J��Z}����gZA��}j^�����Df����� ^s�(�C��[���������,��7/bOW�/`�ɕ���Bf�L����,��ێpY���0���>a��)0�_"��u-0���<g'�wW�tY�&�r!�Z���,���h��M=;7��;�@���Q�`�=���o�1�q�4��p���|���KR��5m$봜%x�(bv��+����!q��N�(�f`�J]q��������"5k〙�%*��!��g�Zd�=�]�����;��x�߫��pC��������|��T�����-�T���f7���9����+o�'z�q�i@���M��s���B�+-��:��p����k�`������vta�����;��oK��]~t&{�8�!&�����M� �'/��}�rF�EC~�Znϫ��"?�TH�Q����Xˢ��G�������������9ً�.��6���aeB��C����O ���G�-�W�݌���]�7#�Q��3jai��!����V�Ն.J¶g���G�Q�C����k�]�C;��f���K{�E��x��t,`�8�{��[��������3��E!8�4M���}�ztߠ�x��[̀36� l<�V�3��H�*VB9��շ]��c��yտ�����#@��y*�vY����7�YT<ooe�)Yi��-;���YXО�y���WgIiiO2���
��γ���n���8�ˎG��q� =���#Z2��<xkP\mu��r�+����M�E���!!Ab#�Dq�2JE7�ױ��kR^�#��&7��D7vwΕ`�䫼TcQ�M�Ǡi0�jH�+=4V�G�D(��<��i��@����<�>���2�P��[�lM�_�����E��J	a���1����Wy�t'�Нε�J��4l:~"�h�'޳�(S�CVu}p�"_#I�̾�|l�jt�#�Aa�zz }:Dsp��H�2�)P���Ď�w� x-%Ϭ��i�k"�	��?��
����$�i7�s<ZHX;�s�>�vcsޕ�������)�T"s�",V��~K��*]����Xk��� /�J��.W��,����݅ӫ��~U.|O�:U?]L���98֜�j�X��,����C��;�����o�c��%���2o �U���<��6�V������U�}Ie�,���W+�%43:�	Gɼm�:�` o�M�>��@!^^ �;0ף}-�*9��5*��(H^Q7��S�L�K�ҋ����<�2Ex��п���@�s%��K�_I�c����:ݩ��'�2������[�»�)�9f����&�y�]��g}k�JD#�'B���h�:�`��T^�w4�s
s����ԗ�����.�,<"��.%=��U֠�S�Y�<�(��&ps�=���λ�+�nx�f>�*�8�*�R�Ұ`4�/hߢiQ[n��-56��p���������m����~{��j=�!6�������f�rUZj�6�O�션�{+"�o���@0ˍ�?�P���5�K6w�H�.2�L���I�1s��'2.�H@��Pv�-6���`����ˁɸ3�_��+I�P�u.3!��;^�f����(%�4d:�[:�%1")�6���B��1����{`�{�P��p�Ai�x2m�J�j�"���x���+����AY:�������?̼eP]�-4�����n���]��www�\���\?�������US5]=ӧ�ٺ��szz�F�.<)M��a�K/ ל��rc�?]@SȬ �}���Id0��ʢ�ʂV.�7%�Fw��E~BTn�Ȩe*ur�Z���t=b���5���z!�s���
��9O.yX�_('%�Ml��ʭTt^TgD�k�Hz�Jy����D����f�/�(VC-�X�2�~i�C���%��8����#uw�V,��{޼>`�-�ޥԝ�a*|���ȸbK����#�lB@XYΆ]�y������7w0�c4N�h; ;*	��R��4� &d�#�'Y"�B��.`����R-���3��b��Ä]%3_a���J*_[o4=?�&�(��
��K�������!���F A��A�_W�\��H����<%���z�v�����(#-B#��_��)�ϯ 5v�ΐ���Z(.�'�}=`v�E���� (٥F#���f�Q_[��Sc�ؚ���Q4W�Ȇ�6 �v��:�/(�#�&����j'���B�i��F�*<���"=��>�n�E�dh�ŮdQk.�aN.�KБ��\�����跌��<���K ���"X"â���/�諷��hV�����Zs_,�6}�{�]�-/�!1Xzߕ��p7���2&�LU��)�Iz}Li ��9�4�G��i�2���I�}/���
1p�	�e�5�h�cvL�,�5���C%C^��v��Bf�Ö3OR�e�B�]'x\w���\&��yO����O���hK������zQ$"�n��)�1�3�0\7I}�N����G=�:���T	"m��ϩǾg�֫�W�o���� �(g� �����~��DBb�N��=]�T�3b�����{5{��>T�pЩ:^�E`�T��[%%8@��ޏ����^��F�x�a�ǥ����E�pC9A3r�ea�Lq�O�#E55�`b��U RN_���ū�}�P�c�&^��"�֫���Et:�brig'?s*>&&&�0�P�/���1D
�-�JAp0c%Ko�y��ѯ���L���'n)�v��r�a,b���h�C-@���aH��1��z/�Ŋ�O끁��P۔Җ��ëB]4}Բ'\�KX����Tͧ�ι�i���~�N}V���`lJ��
��ڍ�j쎕sP�#�40���
�a'h������Y�KRNH8��C�v����b[��}"�q�S�%�D}b{��B�U����_��`F"�?=%�zX?��l�U:��I�U'B��ৃE>da!�"�V1�9Å�6m�d�s�a���R"�}A$8��1�u�=M�~��E�	 �~%��R����RE��*�d�Ĳ��Yi(e@�Ӵ�x���t���Uev���jhD�*�<N\��2�z��f�尭̀�ЕwY�j�Q�S�k�,��<)��������!��������c+a��W��0D1�F����M\@�����%�j�&������Q�؜}/�����HD3��F��㬦�J�!���	>�򋧥l�.�i��b[X|�b��e'��E����c,~��ZH����ki�������u]W��N�Rt��!���lm�)��⼥p�/��\	��#���|Y	��ڳ�h������i�ZlRa����c�Rjrs��� &w�kȿS�ςF�~��֏u�t���a�@�C�@�lDM����A��������K�'��?�-��
��{�++A�'��h/$�Yh��a�>4��D�V��������� �*�nc;*eBw-Ri}��d�$�k��G��Ȃe�����X(
LUcg��n�l��>l����w�7�w�<����{<n�<	����}�{#���D�����4���@g��;k�L��t5�p�̟F-ri�xu_��VS�х��k�e2��Kn	4�Ӽ������P-�80d	�A3���i	�������C���(�����%;���'LO���vd68��_loah���Ap�x�t����Op��������Nf�'�n�TS�5�p0��0�hC���`g�̥3�1��s%NN�J�t71		��#�x{�f���9�-�{Z\e�S�L�q�)��3��-R��
��K����:-cn��������RM=�m�*�թ�șl����s�@�b9p�ŗ���:8a��'xb�g���h�H��&�����j�����������-om�ن�IB��W¦�>$����F	^�Q���MC2�!�Ũ���N� �ћk�$k5��1��F�7�=�.�Z�K~p`���F�Gj����9�6u84t?���Ox\�`��M9��H���Yg��}j\c�'Rk�6�������!��W>䕿/��5eF���pTS�94i����:%�P�/�\��}?H;@qi�3�Y*�~�B� �\���yW�g��G[����*w���b�.ŗ�;�؟��o��ˮ����\o��<���Nw����v���Д���k�m����ھ|�� ���9�������,@h�#l�~\�j��G���Eڲ\?,E�	g�z���j�,CU��c��v__�wi��*���_ؕ�����M��B�;�0wV��#����)a�i��}P�q�^�;�*09��|����Q5;�9���y�K��B�zW�E/�>��K���e�Y��Nʥ�hggGMO�����k�=��k2-�{_NT���vMy�����kZ.�ҩ`q4k�8c����)�ZB��S��w���8Xb���[:����u �L�Tuz��ɸ�SK�*V7nhte�BS�%%M-�^3�V���5ۨ$A�X��&O7G}g33��E�}��222?���P.0U����Y�T�K�� >3�u��c$��-��T+j����\�1��La�-͜���������%S��s���LE�;}���:�t6�&�`�4�{�$�s'���s0G)t���Ů�%>������v7��;�	�+nzv�J���m��-=��()99Lp�� �,��(e��P�!����,��A'�0U��k�k�nK�B�d��{K��D\����C�����3YY�@(45���vg�!dl�,K����`:4;�ڵU#vq�d�/�� 팱�ፅG�#b�h�I\���N.S��B�^�#��ls��i+��a����wr�T
ף��us!�j�����P������<l㋍M%�����7��[iؙl=M�-��� r����|��v����H�?�~ZML�&tZ;�[ά/QL1`�.�>�V�ٹ�jui��۱��5���^�Ze����S�l��#z���𘹑�:c��)���29�?�Ά+^��X���"�2Y�)x"��޺���������{b�����f��)�@P>���9�A��7s(���Q��[X�o�s{s�"�Vn�:MI�W�m`i?�!yq�x5�צ6�茥�_lS"B�sr��+"0�4�Z��}ó�'y�1v��k������o�p�\��rI�H�z�etY�ۻC�U�7�䓍�SP���V#%��zT�4�M@�8_q6�+��j�Ǜ}:D/|�K���l+�"�!)%���ibb�^xz�5����'7X���'��6�E�_���9��u�Z���5����wD�,\�BK��z�+���;bv{��@��	�e�Xe��'�ѡ�ŝdR�}@�ߌ�k�Ғ�m�6"]�5�p{�hm\eaf���W<kyr����dG�����yL�=�j�`�����V�`tO��={C��f2�(��a,�b~0��;��w	u�wk�ԍ$i$��$eL2�2�}]h����i���G{7��x��c-�yFi���aRE+�$=��W���+��-K�t:b_L��ʁ))��p�h�b�8͎���dՋ�b~y���&	������-�{��4��Ѧ����ͽkTw�p�,6�+���aB��fλ��-�:�8�i�+:�7(�%2���L���:�����sq�M6� 	�-��K/����w����ְ<�{5Za]�L��Ĩ4��ˊ7HM�8L��0h����-�y�}�l�hD.Սb*`@R�B�]�.���j�yu"Q�X��RX���f��A�ʹ����.ռ1����:3��a��:V��trq�I"؇��o`;�%�ٴN"w�� V'���[�R�f���kH��sï�FH%6��9�"�L�Ͷ���$^���{�� �A8P�AS�f����v���czv�d.�H��|�c��r�]݈�j3���9�1z}q�)�Ml��=�����kA[���f��F(���������+ZN������4D׸��e|0�]02,v��f���*��v�~��|�,�WrAA�o�%*��wR�+�e��k*���s�F2W��db�Na����"bSJ����n��Ϛ$���~a�X���{]l�'�;��#�2����T`��mi���<~����F�)��X[��Y�:d�Ȱ'��A��^�Q�Z�i�101�A7A���D�X��
��v���,=�7gQ��4k����<��Mz�I��Q��(��j;���WĐ�T������V���w,̕�tΑ�T��x�&��/�>%G���YE�g�n�_�N ��u�)ǝ��-�J�!7WDP�H:�!m��C/�Aۨ����mN��qBp0�\���a��C��H�2��c��������X8!JÊJ�P���W��֤��J�hS�]9�12 ����PŨc��S�O�)� I}Y�T;4Rk��'4^ʶ�a�vǧe,n�ժL�L���θ��:���mEi�G�3��_2F b�7��C���E�����6#l�\e�TSΰ�d`������) Cp�Գ���=.Fp���zI�.�]��<Κ�@J9i8/~��������5�풲ʒ\MWf^�X��c~ױ����� ����+���`ӵ#�C� ��L ���Gh��X�pz膤�"3�������*�)���Țg�/�&�R��&-��0��$�;(AT�����!��x�%e,|�C ϶qn���.�:�!=�oz{{;�ɜ����7��I37{�j8,=t����,t�
��	<��n=�:�4D��j�H�k?�G�&�<���-aqB��g��\w��&
�֮F��N�D��h	�/e1�����Ke���؊�{<���eH�T1Ě�ZK"�i���W
jЯz��eP��/����-����o��{�&e��Az�X���N�~����Q�o\�2w%�P���È��,��*�b_Lx&	�a�9T�v8ߓ]e#c0�P��0�Ӷ��s ���޴ST�y�f��xD~F/��Bbjj�N��}�U����E8ѭ��7Gs�u?����8v��XxX�l,�z��D��}�vF6Ч���9����G#a�_�/���_] [��Wd�c}x�8=�V,ϳ�x��TmaZ���ʵTȄi���(�X�8y����a��^g3+ �BEo4f�Jp�H���Wb$��I([����Ԓ�ꡏ��߰�Ο�t����g� � c6r�/�=Ruba��!G_����rb���$��q�I���F�����7�Ks�𒓓��PlͬhN#h�&�X �t��/ߘ
J�3�����χ*�IŪ��QI� �����Ju��90(�͝��*@f��1�+�Xp��L����� �#n�eDUX�f���qu���|M��c��b�:��U���]���+��*W��@�EM7�3n���4����7_����3d��b$��!���Ґo���{��A���I�9s��Z&C���Jq�����+Ӟ��%!J��վ�!�jܮ����莾��4��:#�"������V\tGc�|�9��w������v�J�Sa��$����9�Q��3(��蘓d�7��k���+�>҅'���O|!R��E�(�Lf�O
v��}D�xz�x<4p}*�g� ����}5�r��
Y�g;�)�*�=��`������kﻘ�N�;?�S��X���J|
����/����x2�,V�@DP�W�q���mg�����1S�`��3�:��cpt~��:���4W�R���<�;��W��'�n����?�RQI�a(��$�S�@���@@��w׼ꈽ�T"�E�j�xk$��Ţ?q�q�C����Z~����a�AZ�y�����@����5�ޜD�T�^/����%=���F��(g��Q�mKE~U^i�=j���p��k��y*E.r1r�Um��� ��U�8�=V�$��#������U��4 {��2��jGS�A�#���p�H漣�����q7ʨ%�.>��/���7��eSQV��E޺&^i�D�˸��t [�#"}��ދ�GR�'�1@@/�*�0�8�� �^Y���y�d���Jc"��ί�n����ۊL8�S�i���t)�?8�L`3c���h�����"��hu�$`�zgfF���a�H��c���J�Z��1YG���	�x�=z��˒c���Y�`2�T�ӒW��A;;)�e�OGLD�,=������O�R�no��$�������)�-�jd6,�7���������{4��d>��䐊1/!۞�4���}ϻ/���X�2&���|ǃԍ�������W���}���?Ƽ�h�����TSc(5~T�	J�#u��Ȏ�D�ImJ�)���V�@�Vc�p��@�UD�r���վ+�RR�Iל��{�������0#��[�nX]	��/�|v�h6��ҶK�F������vH��s�|����_�2J�Gqzz:,�8./���"B}��^��7��I�̛���"�pKNO�����7Bǰ?yo���7+���Q�A��m?�o��Y
�+�|W�xB(*�©�ՒJgGTb��0p�]tc����Q��̂V�L�R��^�w[��a �R�@y�2���8��D�ܤ��$�Y�2��UԼ��	.^�BAS��o����`=������J��r���������0�:��~�B"�l��ͧŖ��H&�92� ~���#��m���#���m�<#^�u�L�r���5�FH�'����*�?�	t���j�ށn-A��֔�7�I�]�(&K����O�jT�XTjo�������y��$$�Y|�k�z�멜�� ��J�KB�Q: 3��J.g�b�qX$O1��Wg�vV�`�)i���ҏ����3%9���C��-��0q���vF���1\�^�p���_���m�^/���i��y��0�ԛ�mmZ����LǷ����}��z?XޘV�wdMmT�Uh�t+W�V~a:a�j
19;;B|LxXT��eYA�R:����Tt�By��Z�*�Q{�rT;�Ƽ>��\����� �D�>7w?��
U�M������^ތ(�쾔�ؗ1e&XZgs���3�Z��jun��
|�B�xy4F���@�%շV%X����bhy ���=_ӫ=[B�^<à��5:)��	�~� �/�z>�hcg��WXX(
�����9�]��@r����y�a�T�AJ�}�9����6�� �tܾO�)Q,�6�(h�ufQ�bHS�"4���aY�`�{R����ښ(�����i��-ˇH676}k�+�>�_q����]�8m�*>]sI{dY]�IC���u���� �gb�@zn[�9"rr�0�h�ۻ\�����.i�8����d:��EL2��֐H7\?�)���ӫx�\�5�U�,�����\�PCII�;��S,ӡy��(��JG�F�����v��Ugu=H9��j&����U}��gF�;	3�B�vj�0?��iww7���oG��j����xg(�9 ,&�H�(�D��ħm�:�R��~����&�����N"��#�F�2�`��Fv��b-��3�oNu�i�}cC��B��aTl�&��%���8t��Н�I�DQy���GTħb�&�^]̲Ա���333}ώ�g-&d"��O�d����a�h�7��3S�*�����+q�.D`��O��.0�>�+����3G�L�1��օ��/�N��6�l��ŷ'��a�
�,�����0+.��D-��[�����j <BリS۾��472I)K|�>7!��4&s�	�/���t���.���!p��c�B���z�7]�JMO���l z*�Kn�l��$�I�����G��ő܉��s�d� 1�6F�t�V,�]�ь	 I�'4fp��՞9c�Kz�t�i�����"�e��unw]Tw��q���`'^�O�)�[�=����:Ȝe\S<0�stG�8�VQ���J>�G�h�ׇK�x�8a�^a!302�H�'i#�>��ྮ�\F<XeOC/X\؜����o�NԂV����R����~�q���ŕ���л�i��-!�(�r�c�a_ey������W@յ������+��Pϐ�Ɵz�3[�|��Yps޾��ʗw�x���Mľj���~�Z���&�t��"�T.X(�ȍ�>M""P�5��I�S����x�%	��ib�:	��Aw�q���h���F���:��ೌ��b>kl�j��tm1�v*��C�U���^���G�'I4��1���t�d�հ�=��[q�j���ʜ�z��+���؉���Yb�P'��[(���h����%��O>�,'C虥��0<��sǈI�Dx( ��E���� =	7���R 1��(:��f���,o�F�_�O<D�P������݋��]�� ��ը���_�̇��b\ŝ�0љ�u���EL�e1�9�4��~�1�I�ݩ��%�cNO�%����
��9t�s�$5�!!%?�bF��,�B�`+��b�H*q-�7[K,������QX�w��86k
����]Ƥ���fie��	8& sP�����3��-��I[���+^���SC"�օVRO5ǽ���8��w�� ��$Cǜ�Ѽ�����9A���bc�@HhOVn��4�о��0����]�V��gR�<��0��2�'?j*M��p�T�ʏ�'��YG-sNb���|�.R�����Z�(��.�e�,q���$;����ds]��]򲾐2����:��!.e�1
om)־{A�0a�`�k� ���ފM����<1�#{9�ˬ�X��Zm�`�������q�`i�g�M���-��q�%����C��&��t��&�n�AF�hT֙���|����d,��	���4r��, }I�Fj��;vB�
>[ô���s�fY�#���E��f��3�����`�q��O��:�Ȅ:��[��݅��i�ǣLts��C���?����:������)"}�:y����j��X�r�����O8�EEQ͸������7�2�)䔡��|v�4��!�]n�F�z�*,��a��n�X3z��-������ch�Wq�沄����<o�,�q�ߙ/���;���>�5�������qC��O���b�!y��K��45a��~���"��Ǐ�gWy���b��1 �_�&�t�2?F��i�����v���a(��گ*UN�pG�����C��>�,�_C���U�_]�H�b�1�߉�v������X������A��	��+
�k}ݲ։�U����{��l#�!��d��3����1d�'��҅p��7��/��!�S�G1�(�V������bɠ�H�8��*���x����	gx�+�%����0AD�+�'�[]�Rm�JE���t���4���=%�X�8@m���VN��Yu��C�m7|R������Y�O=]5X�*��� _Ո�	u�-^ǋ�N��J�$�J��� q��(>�k; ��(vO=��sz������^�d� ��T��LƟ.���o�L�k������B�j�C���Օ�ʔ��`�HX��K6簏�l�³��/�����P$ �Q��gXs�mWy�p���an��{6�	$���J'��P�t�D�	f�pk�d
���!yZ�ǀ�+�ޮ�J��Vǡ/��/�G�.I2��Ƈ�nJ��N��jWgA
|ƵM�Ex�d`T�#fM��t���{r�<��$)��"�Mia>���Ƒ�,���$�}m _E�yn�o -I�Ut��va��Hx$��)���JH2�m���:�4�Y���(�L_?�`3іL,@�:y`�g�ͷ�Gi��3���z�џ>�[��-�/�^A7����������"���-b�d�m�����w�>�Ҫ�w\g��ܶ^������HR��{�r�Ff��Z:�#�^�N�
w�jb�\�dBm����9E��o����L��
S���2 �$�VC�n��<����%TȊ�~v���@���Cű�
���?M9���$���`l�`\i��Pv\���� +�Wj;3��y�<��<U����aC��C�z��P"��R�
����/��c(V� ��(��7�Ǐ�K�NkU�ަ��P_���3��o1m��}�jxf+��M��s<�i�tt?#,�s._6�)'M��I��L\�:�őC����4v�4F��	�Q�sZ��Y��ۅ�_�=�9�9(�	��E5J�(DtS0\2P�P'�Md�/���\�OP6mj��ʄ:�`<�X�z�'R��э35�)�U�⩹�jNv)`��/�y�\�{���6mM5/�b�@��^�.�	lܾ�9�l���\\� �Ux�,dם+oa���H&�1��WꭴA�%�Ř���b�S�oǺ&���J"�;b��h��+1/ 0�J��GqfB����RM���!�˘��m��x���J��$��ZΥ㢶>�@�1�	R	y�&BGĞY����m��8� �D?,R?L7�����"�,:�(�F��9ܸ-���7�|����Y�p�ߞКe�:,��_�!Q�H�~����Afb�%D5��_H��,�ϖK��WkQ���fG%a�,�ef�Q�����d5A�^<���Q����ԥȊ�	C��X.���I�Q�
\ΤH�L���Ф�2�ʸǩ��e�_3��To�&�[9��jة��xH���h��P{4��~glv��r�ƛ�ܞ,٫�%k<���0Jvf��>�[��o,�"Q��ڶ�����*�H�	�kP��0 ���2�K����BRŞŝ*����$��J���������9� �ە��Q��\"c���"����>��'����+��xe���ŵ�҇��QM�p�6��!Ǵ@*W/⠧]"���'֔�h(���ֿ@�f��`���`j�%g��/8�:�^m�嗟��B&��[q6����5q��z��!��*��<�z=߿{=).s����P�S��<ʗ�O�<7(��/�)x ��m���\ ��k���4hݯi_7�yW#�j���6��R��C%��M��xO�$Ә��q[�������V��v�
����N�l!��Ls���RZˮ����W\���Ze��[%�3%']u���Ԧ�xz}�g�¨�=���`���}x%��p|J�(��.n-���{���^~W1��+��iQ;K0>���s��ye#]1�����)����4��90d�\����pNr4�yw��Ѿ�]o�k�d�
���m��_�?`:_.,��h��	���u;I	*��k>��΢*��B�F��S�7�q6 T�>c7�R���K|�/��sU�����$i[������o������jϝ���Y]��Sg�³�_������C�W�	�㌏r<؆��UF�<� ��v�r�e�����W�>�:_�yꮎ}��l"���Q��aD�BԞĦ��y��N�=���7��+��:�|/���8� ��{���LJ���g�9�:�g��b��RbNڛ�O��TK��F�F�+5��׳Y����qT�Ԥ	)Za�OkW+�=��	T�|�\�(��m=����hM��Bz�yb���"�w��2rc4�|��sﴙ��V`Dz/�.�qA�/�Q���+�̼�P��=*�(0+�-O�+�%����n����b������ԁe�E�e_U�Qp���јZ��rL��/���8����`�]a����P�H��ɳ���"ȗ���+SWs�}�i���sǥmٖ���=���:���+�!���nv���*�f����ԟ޼{�6�>{D�imR�1~n[=nG�̥W�/�/֣)��<3T�G���$�0I#� �'��pE��ki��r\(��.��{�<K!UD[?S:A���{V/q_ӑ����gI�~Ji%�WMJ������:��	�1|�А�Z��l���P�ǵ��Qᵦ<S\ퟓsq�>��K����X+�m�Τ=��.A������)?������L��.Ы�`h���q�)-vHf�lg�Z���1"+N��������ف��Iͧp����L���E"��6F�ҰoZv��oJ��QL��J�n�v��{o���bkݚ����� �>����G�ҝRW��a(T(����405�V��qXZ�)�S�2ͥ,B�L��Ha|����Z�gٸr�H�/���8�Vӎ/���lacs�L����s�{�ړ[����ࠫ�[������:ź��I�-ʽOߍ��%�s��@�SW΁�`oG�n�钨(��k�#�G���U��`8�`�jx��r<Ý���&�`)۴ <t���,ŉO��E�=�jd}b}��|�d	˥����G_�9O$��nE��dH;�<�_s���X��	������)�����)l���ja���QP�HT�Ą���K|4�y_'���e3�����B^48P"x�b�twmYu��W�{n:��z��3«/q�W��W���^u��y��devg��-��+2A��nw'�l�i��A��@�J�/�Y��s�AIյA�(��r�7R�9�_�#u�E|�vZ=�S��ݘ��!Y����z�S�=�kL�Xy�Lawq��a�>���;���I@���o��R�?�7�,8�,m��1�x���<�A@��_vLk'!��ԈcPMf�CB�u�S����@ۜwW�};`qFz^U�.8���7�����&I<��ٰ�Kx�����?�,~5X�w��q���b�z�W��z%mЮ�>Ȋ"-§0ߋ,U�L%��>l�nӲj˙���Uze=�d-Y&�όQ�h,������ 
mgQ�S>ە��voӯW�jsu)��`C366�K�F�i��:��х:��ک�Pvn�Mͅ��roP��$ ˀ���!�3�1D�p�߯W%�,���T���;$��7�=�UL�HU�æO�G��i�4lZ��:��Mk��EI��Wsx[�S�F����+ʿ��
^[6|�N�4ʥ���1�͊Lj�'Q��d �~-�!*�-XA�E�N�`	$�_\Q�:�z���Jx�u�*��'n��7HaJ}��D���Katq!xe�5��!:wgi���kߦ$�=/)*�,'|]&�;�%}�I4o�t������*�.rv�$�PcK(� e�i~&�V���\(~�f�ZP���|���Æ�S��}}U�JZ����#OG���Β���DA�k�Vj\��5\�h0(aSҪ
4�����@!w��~�;A��MOZ3�M�&5`O!�������Dά����1m����d-KEy@�_0܊,v1lG�J�`�T����?�G�������/mHM[5 9:[�%9&��?u᧚�	=��w2�@�t�aʰy;ɖ*��"��l�u��עs.-���ߓ���Ҡ�]	L�M�S̐1�Z`zc�<R�|���Nz�/�J�2[���)@t���<(h���|�RC#Q�Q�=I��� x������О�
�{��!z��.��[�������z,�é�}��YT:C6u �p )�ϓ�y	`%?��T��\�Py�3�b��m`5:����@W�����O��nH=�v)���N�Ɨ�\;��6�p&�8{�u��Β����+�i�E��g;%.�r��;XC�}{�� �ɞB#l����� S&)咂�����j�mH]�~������e��'��|�6WK*V��٦�3����j�pR��%c�R3��c��������ƯD��b�	Q�h]BԸTi�Q���K!���r�;{K͖������dlCbt�w�wu���dxB�ZU�C�0u�`�NLX�q�3KU�JJ�@"�/E�胃��ꉣ݈g��s̙v�&�:��94��r�>'2�W�_PM8#jh�z���_\vv�>�����I�@U"�>Bx�L��Y�F#��4`2E�OpS2�\����j8��d%�:z�3�QC���0D�p�bWBƖ�A��ՙy+q�����5M��H�.���^]�r4����q��ӉF]էit�b��V3e�p��R�tE���,&��
�܈�Eǭ��Z�yC��}t~	���\�R�� ���
/����hq35�a�?��q2m��}Z��ܨ67�4�D�[�1HѰ75�j��+l�ڪ'�@��t�+����-��},w��ܘ��%�#@9�fxkb����ih���,�4$��#S���������Ueճf�*/�u ���]�=��1'��<w�C�{v$@
���rY�� @ �TZ_�ѝl,��xG�e�%���{���!C�lך=�&�7s��㓁�}ס����.�>�6�8��ƃ��6�����@��4Ҩ����B�>�T�g�w\�@\�F�yL߇�U~�M`g���ڬ��ݧ��!n�Cq�_ɝ�����QXq\ 'Q�YFJQB�U#�u$n���1��a6��5�gB<tvT�f����FX�E�4��>޳1^�U�߸�J�q�&�U_�����'�,x�g��yHw��X|���͋��iҥb�.�"Gz6�	S�4z��M���������^p�g����Q��	�6�{[�r�t �m@�釭�G9S���;D�r�	�M�uC�'S	�FB`��v7�����i}y��܏��c��{�>�����v��}��׆ݜ�Դ,��?f� _�ˇ�e�0�ȃ	;�}�/f�����?��4G~�������#1@��;�~K�W�����B��A�v��苮n̏�]�e�$������[xt����h�%'@>mʽ�y.5�H�a5���7���O�CӶ�%�5wj2`'U�N�H�	�P�(����7����	���OVN4�w�ɂ8m#���L0�J�����ͽţ7	D���75dW��E���ߝ@���m��όuH������"	I�l w7-ll�á�Yeo�$h��S>��6?N��0�xԩs&8��o�Uq3�:���1���� ��2TXS����sj�~axR� q���[�����P5ŷ����=�RAj���u��~�l+�P�9xVU�,�Y�i�h*f��l���އA��-�&�#�k~Mx�A�E��ؕ�I��RW�϶��s_P�w\_+���U��𤣓��+%z�	�9�~�b�����]�<�Y����R�<Hy�s4@0g_�i�t�(���XY�zC.}�r�B����}����/��ő)AR���[U�H�j���Jhh�R�U����5����ݕ�%��Nn�xD�6��[���i�K����Ga�Q���=��~Woy�l{ٱD��[�/:��ήE�J�nܜ���g���{��b��Ef�f![ $̂j�of2�o|�Mmh�V��d49�i�$��q�����9�Y-6��咒EWy+/�>"*�r7��R������(<�m�є<еM����D��T�Bu=^g��>�W�ݒ���$���8/	��a�5��;��(�~�Q��8��.���P��9`��J�����EK��0e�Wffv�,�R~��JLT!�%4�7�̌ɿy����6R��c��S,g	���d�����W隺o5V:b�}3���6rmkhK���/H%�T�qe�1g�=�9�Ő��)��k�V��Z\�WO�JmW2l��O�4�)/�ݼ�)�$ѐgHE����1�kO���W�抿9-,e)�d�������.�Zq�te�J��m>whՈF� �E��h43VC9ǜ�3͔\�b;�7�9�NG�t�bhmnZa�Jy��Z䵵5Tt��
&��*U��T1��J��U�cQ�G6�3e*vt3�DŤ}�����i($���K�G�#\ӄ���c�r�\Hɓs����
;!����������	��w��.���E�1Ŀĵ�=�:Q[n�|P�ҝ{��?&|�+�?ư�	���SH9Iu�A�nn���|���T�Rb�O
:֢3"��D�� f ���Z�,B}�]UHga�j������0R(��Ae��p��ϩ�W��=C�9��a�83ĵ+]>�X�LD��a�9��i�/�7�=\7��IٸH���=�%"uBӘ��~��	 P0n��3_�7�}�Bqiqw���Zܽ�����Cqw��@qgp-�n�=����O^�JΕ����k��dFp�XfddD��]M���t�7]h��Ҍ������B�x"	��Cq)�D$e�@}
�gA�Pe��_i��t���*)#�2q�݅�^��.{=_���O�Ff��������ϫ�a���p%wʇ�\�	-�$FW�H�H:T��m;�D��H6Y'�~�s�l���>xݲ���H?��	,�pmxܤ�ש���Ef�����u��+-�<�"�o>�}�[M�"��o��J��0{�<|��R;1�hz�% q;��2BS�,��]�j�#L�8�r<XpӋ_�=e�s���ޔ��{)��ڊΫ���SuJ���#B�<)������@z�Q�I4i1��c������<��Zq���6�Z���޻������}Y�Z�!��+��WkT�à:�����(�И�����Yh����9X��)�{q����G�7��xæp���a7׳�:�����&�3&����S�m��|��
�Qr���ت��Д��	�}�ӧ���D��r���ܖ�-�ڈ�*0�ܭ�ƨ�p@9�rw��pD�����9*��^�[��O����X~F
97b��<��2<ײpss���_�kf'TS��H�e��G�x���}�{�x�Z��{�0ϻ� ��HW�/�	jX}a�ٻuk��$�/�W�i=�9�+f���"��ҵ�AT���.�VV��hoO���}
���T��1kY�^�w����|�8o�0"rRRRr���vW}$���iM�%б�g�_�����j�ƹ��e��z�;M���/ٲ���t9q���2��Dk�ޛ�Z�2������X�3��jS�zU�NY�ˁm,�����L�Yl�����"m.[�tDd�JS�4��uK<�hɺZOrb�Ϸ�1R�Rc,���̊���Ԭ}|R�3<#������g�ȝ����q�x�).��([����",����ٶ��Z<�Z.ؤ��삒qm���v.F�E�]���rj~)�k��O�F�χ�V]��q�����?ֲi�zρs��0��vj�W�SP[��ۚ1�{��%F��au��&!��9O��j���JV5t�(�
�mi�]v;�K�l�je����ZK���.�VWNS�s��Y�S��+�_��;��.��gq��\v�z�~�o��%!��g=ߔxY��2m�&�R\|e��7�f��3X>�
N>��uQJ�ð����C��U%V�^��׫����R(q;zLqI��)P�p���>3r�J�	�id��r/rϳ�\J(��A�1�v{.���	�%�/g=�b�o%�veHG"b�/;D��5&wg����q3b�)�v
�G���t%��gzy���Sh����<�I{'c���a%����x����f5��I*)��U�T�{���B�F򙗖��c��2$�6p�6A��o4�ʯ���@k	�<\1�&L�F��7��֨��X���٦�,7"�n��kmB�Q8{�ҝu?S����LkCV$�78�O'ԙ*2u�p���I�Uй�7�d�͹v�포R�����X�o��˧"N_�=�2=��֪_X6dD��n�'2ܡl�QnF��!+�@J���g�Rqw]ܽ�Xry|AUv{�8r�yYiOm����W��x���~�/ګ�}�,�Nt��5�@�_Ț��/m�y�o�2�3]��WV����w�[�ꂀn��p��"{I�|N���%�$�d��}� �$������yIΊԺ;������q�{��<g�Y��߈O<��n勭hZ"�j�Y�K�UZ�)�(�"�\=�+�e�"��GD0�_�E�ߣ ��^�Ɠk1�Y���ɗ�興j4�7(�%�{ZWӝM�s��ױZ+��� ��\®�Y5��[�����m�z��b����L�Y�׈>˵J�qv���j�rWM��W��xf�[�O��H�b2�v(1���e)��._N����Y�C��s*��m�R�%Z����5!_�|6UCPT�qX�HH4aރ�|��JW���#ܹ��^��3P��n���K����kB���}.��f�΂,���������H��Ŷ�@�A�S���X��t|�ER/V<�s[x�4�:nu#|���85cv`Ԩ,�<s҄l0T�����.�S7�ч�@I��S��2�żs(g��b��4 �lH?#+��@|W)X��4z��W�;*�oC �Pv��ߜ��o��y���5Ͼ�/�h��רI�04q��,���G_���n
p���9/K�66�\q���yA�&̖��Z��<��[h�<�/B��._��<k[��w5&���J='��ۨ+NvҔ}*��mJ�D����A�E�j(�P$$�3��݋�����?�cs���L��"+��^�[-���kM=&���?ɹ�H�-{�[�����׏L~MJ\�@]S��X��T��\�a���&���j+x+Cɲ����Zޖ��5ed^�l�>�pDrJ�h��������IԂ:�(��Oe��~�+�F����F�����E[[��?��+O�C�2:,{w�2��d -��z��ǳ��.��X�����n��x%ˊ�� ^� ��GI���1]y���3��+OoǿW/\�.d7�e�~�c�k��c4���Y�:�q���|����WJ�\�Ȉ��[����X��OW-�)�ax�S/7�ĕ��wS} U'�,G���}��P�8a�r�ǥ5Wi@�yj�/^�͕���!������p�/r�VO4����>������
I���0����ěN=N�n�}�(��ў��,��L��7��<�������@:�ɠ�ne����T�.@�����h�ͽ��BL����t�o�1[o�4Q	�٨P�P	K�Y�E�OA=�s"t��j�<�a�jbbf�]�+��Yt����;��ӧw?ST�0j��a2�+Ύ�l;�e�L�sU�:.�|����Kt&����vTx��U�y�����8N��i�_��3�sS���ք��H�x�,�c��0�tWc|f��ǃ�z���;��U�[��28����c��<F�4��.����}�Xi:�E!�G�9m[��g�����i����T�+�67����u��?��·�P��q�X�s�\�!gƎ������������h�����B"?�C5����șR<��� ��@Ўvص��ڱURђ�]�%E؆F���Ɵ�\����-v�z���/�i�v�����M}v����e��khҝ��� r�ۯ���D�"jᓒ�ͽ�!��/ǩ$�������<uu����æ|�g3å�d�>��w'�6c��.(]<}��ut��-/RR]�oU3�Z�F3y�9i�/����.eP;,ꤾ;f�"�0c
y����,5=J{�Ģ�н��ֻ�^�����3h@���k�_�9����ȋ沈�
v|}���5=+�dup�s/	�䄶'�;Cq�<�"�w�g@��A~ϳgL˳YOYKr�Z�������i�k�����)~Y3��ǻ��"@�p�)�*X򒲦ݵ����`��Uё~�4�͊Oϑ�#��H�'�������\���oЕ�םg���=��;;r%��=9|;��p����6k�2^ږ8��
�125�ȫC�Ӥ�A��~s�̾?�9�\���9yo��"iI�"$�F�J�[A��M)tk��7�s�
����@��/��Ƶ���A ��������n��^����lQs��:q�)f~�W�����p�[��Ew�c\�j���u!TM�1;����{!3^���{�R�]��2��E �p�r�+��Să~G_��I��ug�Ob��}2>PG��rڛ��6�?>Q�k�9�.� O�/�ɳ��c�@C�K����3�:�.�ܓ�@�u����/ĸ�Ʀ�ً�d[s�c���ԍO���Ρ�U|M�q�U��bYd�4}������|{0���Oo�n/�4~8��z��H�3)�{i�6�I0a���V�x�6�����[NuI�	��F�U���+�	�q��Ԕ?'$j�r��n_�&16M��
AY�,̕*�a��
�N=B�[��x�F^���	z�/�OL"\�2�A����S�J��>Mݿ3��j>Ɋ�lM�S�����vS��:��,��$��H�LH���_��u�X��N��s~rSv#�?�Y��mCHP_������ΐB�b�Ό��矬�ZU&��h8��'��5��\�+=G:�yl�Y����+>��}@�����4[�V�$�/h���!D���#�
��e|����d <�$$���% M���7��pa���Y���T�JTRҨ�/����g�7�%滏� � g���]��ߵM��o4��щ����I��F�!C""b���o��~)�^�[}	Ҁ<�^G�=3�f ���	r�,{���i�S���(ю�T�@j�OMkՌ����5y%����?/Ǩ&-4]}�,]�(o�þ`�hk������̺=�;�`�9G��:����y��UPk��)�s���>&Mr�ٷ��s��0�L�(�����A5R��B&W��^,ӳ�����sh48W�U=�&.U����7�/���%~?�Č#T�w�SƧ�Wu�x/���um���}^r�����j*��©�aux�P���dҀ��nʹ��PF.�Z1�� -�߉��&?��9�i�(H�������j�O��ѩ�UT��j�{ڠ��	F�z8�lo]��6�Y0MѨw�qL��030��	��Ĥ�T��0%�t�7���:��BJ*C
��ߥ�)���:�7$0����	�s�.�FPA���:�eǉ�&@��r�7���A��K����>���X�FZG��?���%0)�O��2�IA���j12�~+7��*'�u��j�Q\��ed۱�_��ZЈ��=��zqm*�5����sJx}X7�!��w@&��Y{�����쯦I��B4����y��Q��0�_���[�|��I#I�������k=[�s����������=���:n4�C�UIԨ��v�����{k���.|lu19��S���^8��;O�N�4梱q<�t� �a��#qc��{��}�gc!�w0�v���\8�d�Q ���D���4�yF�����V.u�׵T�}�0C��G,&����O�A���:]���{������� qB���<U�f4)�ڔ��?�%����<2��8e�"jȣ嬄�8���AF�g�e�|�~�z����!��s�vt��9�o9u��D�+D�A޷C�Z��y�td7�3Ӏ�./�yMu��Nɰ��E��r�����w�mUP+s�&c��	~����vS�i�zt���I3��/��m���&,��:n�ǔ�9>GF�BG�m�_	�"�͹h������Q'���2h�+�`�YҨec�ў���7�WT��{Î�AĢ-�.�\QO2����a��7���P�>�ط�����N�{6ڃ�R�@�����hJs2��R��z�|]���=��$f���置k�1+��"�V�gF�؝E���VC'9���t��OAE?5�fA"N�@�>u���z�T'f(}_N����H:M��-�D�D�|��˟��[��Lh:�3^�S��.2o�B^H&��Ȥ�d�dԢ>�����^�}�����,
E�M�S�]d.��)�>	j�Zb�|�͹���rS.1����xN5�i� g��/��o�l��������N������1}�f�J�Q��D��7�(�i(t���:��x9��sq
��i��R��;f�gE
F�J��,�W3�9���+��H?�7�__���{��ĵ��Pb��H��o�h�Y;i}�@�,�a������|�����MZ�+��Δ��b��z�K�H��f|>[ZA� �����^�V��4"{2pE�<�u���e�ƴ��'�凢\jp0�;E�|��o��琣��i�P��z+�]sp���&vtHl_����V3��3#�	'j�>|�C~�emͷ�F+����_!���y	�.�O��i�Ɗ�o�ڥ�oo��-&`��^�[��x���� {����7�%�ɪ�э.ⷬ�+t�������ꗬ�ɭ�Ha5Ż3�'�R�G0u
!�s�C�(�C6=��٤N�\������Q�^�`�A<u�
?�[����S7:"���[��_O�g��G������[U�Ñ�w_���%��"�֡��H����o.~����9f�)���&��~��t�O��aq�~��u�K�e����BJת� r����=p� �P�Rh��:}E
����~�H>Q ̦�j�b�#v�G�
q���q����q'�_Y��vHlގ��rx�_�Ir7.U`n'M��y2�e��y��z�-%���O/2��x�ޖ[�\s����EJ1����n�n���Xv9Q�#����]�b�VA�����8Se�x���}��?��|9�d��o����tq����静c�N{#�.�+�}��Q�5c'�];5�!t��&I��S��4Y��)gQ��,E��o�`dQk(�i�şڶȺ�'vg׸q��/�e�]@��K�gEP�1�԰���N,�9��k%@@�:��瞌�i���=��&���oA��u*��{>J�'��	fm8�
���W��Dz��^J]ء��y�����f|b�3��fxwP��G�Ӿ���o�O��:�������Y/��E�Je��(�r0�
�ɭ �Z�72����e5WW*
�m��o`⩸O
�J}�g�"|��]����[���%Za�zJ�Q�B��lSf|�>��6X����veV���7,Hz=O�L����&�����[���&?2�f70G��WJ�����Z^n.`�c�@�����������س&o�r�1����ʃ]������aV��~�ovCB���3M��`��(F��,"aѬ�T<�؄BZm�W�ԭ�y4�?I��~���-5�JĲ`�ez+��v�=l�#���3�	�Lʚ h3+1\�f��K0��<��b�h���ML�+�ޔ�֪��x�H�2�]��p�x�"��H�O^�z|�?L��#���j��ۄ6-X���>��m�������.� !����Vʙ���a7��)��?f���%h�B���)!�5�oB������z�{��$�U��ʝ�c$=7����+`�xUn&!;�uJ���᝽��U��1r�i�nɚ��^bU�G���g=����q��n⫟��ܮŞ��u;�R��T������z�og���D��֎�7y�s��l|˛L����߂x�w��N���+ Ϙkf��M��1�&"Q������!P��d��]oKh����$�������B��:b�D�����y��y�N_q�W�Uor��e���;I�����)l����������=V'r�z���G�"-��9�H�����w���!�)*{���P�V�Ŕ���z�"3�v8��}.'@�zixMrJ��Q���40� ]��(}U�[��R�ٲ���{�:_�=�]�w5��/�F28�u!iL��1r��e?t��2X�<���.[Vr"#e��p$�$2wf���갛'���؄Bų۴e��-�$~ˇ莨��Q&�-�F:@g:<��̛-*G���Ӑ�J�N�p_ݳn��Q�mRs^RP�p���X4
�0_0?<�u-�0�_�����z�3�>���vb���u�,s���c�̳gk�jR#[ZR�v�>�duaM�ޕ	����4�d��j=d�c��	]B|��k�-�������b}�ܲ_������}D���%�1�ک���]���C"�K�70����j�)<���Z��.e5H��8Qz/��1R����X\T�k�0r���6��	��Z�ȥn`�		'	��+Q���}r+�j%�A�r�a��g�vx��~]#�J�N�ݤ~; ʲT���|���|�ţv��۹]p͇|�ћ���FS�u��&��cc������*��5:���DW�@��<�V�â�����0���å+��(p�4�N=��b
Rnq��?(��Jv���C�glZg�/�Ëi~V�Bh�` �k�����|_Y�U�S��N���W=Z�{m(�Zr�:�0
�!c�����չT#��>�>�C�{ �_�n�6�-��G�?�
��f���z?�3>����V	�<m#Tԁ�`oIM�9=R���Pw�9�l;u��
������S�-�3�jA˚[��O!� ��ȁrCB�^���`w����~�N�)'�M߷>W~7%3,�sj���RL�b�A��Ft�	E�C|mF��{oI��i�7ڔ��3B_�À��ʸ�Xd����"�"l�����r���HOo�V�DY�}w�#����6�6�N�7ͩ&}-���V1�V��q�Ɵ�֬�(j�����Q���8������si�xl\�4���0=^�U|q{)Vx��3����x����{���%^�]�Z��ݩ�����,I��ǟI�=�UӶǫ0�R]ƽA�'�.|�.�I���=NL5t�~U:c��&	9�3�u��=�>E�QԠ�ssVKP�{X`�uP骽|,F�o� =H��&���>�|P�\����c��pX�p˪.y�s�z��8�)G̻���>4�v΃Y���'�RL<��'q���"ԙش�������m����S;?I�&QR�u9����������fďm-ы�"��B�p�4����[0���w�{M1�񟖖8�O��<FHX����M_����(��P�YBPc�[�a/�1��}k=���\�$��jL���}Udn$����W}Q2��9h
�g���+�#�C�u�N�7:��S��O���hL��2P�9��!�pZ�B�]���)�5yXܓ��bG����6u=�G��Ҷ��5O!�#��H�M�R�J�$�T��r:7z�\�����j�l�T�pu�1�ſ��%�M�wS�e�FBW��+jC1��%���,�u6��Y��7�g�jGf1X�/�C���
^x���6ǎ(/�t�x�]�Č�ҏR� �%>K\VV��K2�ə�J�gg:J�
V("1�i�Z}N3��&DE�)�����4���G�c�<��p�O���,X0�H@̓�����C����	��Tƌ�j��D��	E���
%���b�����J*w�w�}�{����ΔK�z�nxt�o��D�C�"l�#ޭ��3#��v!V�l�s�����!:^�� v7λ�,'?�o��jO>��[|�	�:7ѕ?�M�O	���\�?���J+��ڝ��w�\�}���1Pc9�i���PN��&N��M!�y������pm,���{�ԋ��=?5�(�G��z_�jԿ��FU2����Z� ���C@�;j{}�O�PA��%�l,/�z������+���ܼ�K������x�-	�:��l�4$�bS��G�#N�N�UБ�����B�t4�u��k&ˆ_�TV��8���?-v�}<�2xN��蔧���x����<�ȡq2����b������x/�� �<�,W?�g��/*/�5��m*]�V�J��)A$�{1S��$�
�F��~c>�y-��_2��+M�0��4�'.\>����ŷ��	��6�"\u�nO}n�F�$�}~iݵ!�_�U�t���_�!������g+��g���{(w'���a��.ox?{�O!�K��I���히����h���'W�MYт�p����F�O�#��ʋh���-U��I����RjmSsX�:�Ze����	;X�F�E�4���;��%�H��
�����ғ<�zw�Vi{gG�� $}���}�]_Y���6pc�����s�-M`9�Ek@`=����-�H�P�	*H�f�b*�XT�Z�$�@'��Be�Oh�^ɬ��R
O���H�.6g��#п$�~~)���� @��+j/����M��`��:��>�&�à��gNu�l�ͺ]�p#������ݸ�65N�����1!>?Ʃ_��z���3r�Z	fX�� ����;�y)� ;���E��T�!��Z��q������9�ѥ�[Gք^�'H���N
b��X6L^Cx�L��(�dc���`�,C�Y�M�&##p�2�"�u�"js�q�RuGb��j��eW��C�~n&1�Ԟ1+13��s���pb��oؐՌ�^
��_���X�̂�)J�#��Y|�9�P�"��7�/���	h���:�,��ן_S}�P/�炄70�������3E�?y�|Fm��2�i���Z�\<Tyj=����aA�H4HBY��HzL@>j�8[)�'�ɱ�#��P�S�ÕF��y��:B�2������)�5�����`ɞ�on�F�f� �d�N߭���BY�{/�b�m�.lE�R�:��}3 �J2⡜�R{]�ȑM/*WJWm*[��(���z����$K�q!��}������kv��7�v=my���n>/��z�[�@!��-��U��_8�qo���i�p2�$���%�N�����pĄ�L�^��U���m�d�Ѕ^�@B^��d�vC�����=6q� �HO�ЧGޥ��:� {�Ƽ-�ob�����%	��ڛ�Jٻ��'߄9�/��>/��>;?����M�fA�9���� 	���O��!��&	6�J�1�'c���h���T�^��"<e�6���������.����ڲ�S��0���{R�: ^܎ܻG�+W��'3�ŷ *��A]��<���^.B{�)A��g�Ō9U��7'v(�r���h�^5ϕ�W\��=ºUH�J�v|�=�9�&r�������Kwt�{�H�����E�&�fG��K���NK_:�N(}� �����x�V���p�ۚձQ �K� /�e�5��V�q�՜�q���b����H��RK�����O�n����Wsyֱ�<bp�R��O��P�eh*���-^cjxQ���J�	M���"||��� g?�F���%���(Zg�_`a|N&��� ��Y�]Ð�m��7aE����|�y ��G��+1T���[@������r�z4t����h�P��u�`x�8y*��]�k��b	����ہ������z����E5��RJG���S�n}3�<e�&�_o�3�M�n9i�-�!�<R:��\�'&T���I3ۢz�f0�d}�	h�;�fPh�"�#�P��(������3�2q�Hd,��6[���P�����m_ƖBvۮ�Yv��{�qМ�X����*�v�CBlw����9U���.�#Cn詹�:Jz���B޺��4[�[�@����J��:k��EJN����&O��1�Q��q�!�I�*��\�F�9������W'�5n={դ����E
U�'�Uv:2Q�&��σ�듊��E4���p��!�Y.��`St�v�����_4�0F��fx��׻�)J���~��D]�_-?W�o_Y4"�G��[�>2��_��y���}_��q�Y�&�sh�QRh� �"Z+�^�9<}�8ŋ�3c�����`�g��6K��O7mw��RyC�+����+�8�T��j��q�|�՗TVs���Ek<�������[d�ر�Iӡ��ޤ�4n$�С�
G�J�EPS@9����;��zXn����<��ܰ���Ќzɝ�1��5�`�������L��6F��X��Z�~��t\~w�3u@]��(��7���H0�P&}��:Jh��+�o�w����:8�D����#��W]#K���y�o��(�JI���}�ȫ�j�B�+��pw �r/�P�$4�呎���_�s���8p�,�&F�*P�E!C"}��
�ja��V�G���\�6C�@���V|E�d��@ق�J��_�*.����s�"m���@����M���2S]e�8x���K�Q��$��qz��(�H,�Q�������
R3xZ�Ogj�R�]�������p�}�Tbo�U ��_�v��Q=���	-�8ol��Z q���ȿd�{7�S�<��u��?;f�����_	�c�P���7�L���@�t ��4|!�\��L[)9�����+�h=��{ӌ�M!fv�:�r)�ڧ�C�:|I��3g�oB#;!�%�f|'( ��õW�l�L(��5��޴PPPH��G��fZ��}�g���Fʨ7��a+�?zDG'�@,Xj��m��g�z2���um�����K PEF�OW�3K�\�=sU�R.�lx�=��:�:|Yǹ�M�����p-s�e��L���n���<���5��csu��_� �����]{����}k-�h������N��}baH���iT�a\������m�T��E/��E@^�#I��W��^����aW.}��+���:�$%�.[#�^�љ#�ٵ��o�-���ّ��) ��-����٨aJ-!��+u�]8٭O���sRr��E� 1�al�	�@g��S���M��R˹��"�#_�{X%]I��h�����"R�	������H�۳�O���	�~պ)F�65>�dU�h%�a(s`K�4Y#ѡ�T~z֟���3;�����Rv���Z%0"w�,)�{�3g�h��E=���g"����!�7��!Pv��H�<k�l4�s8 �0�B��~�U�zzz'B�����.�u���9��K�%&׎P���9��kx{d��&ee�Ҧ�E,>�\`\fz��e�x#�P���Y�C�!),�5,���'6u*Hߖʉ�9(���&"	E�}F��x��/5v������ҹ{�<���� Ŧ��*$,��0eU�U��������%��o_���������ڻ���c4ɬ���Y� !���w5�D*�`Ń�Y˅N��N���*���Gk𑹢")D瞴��#�NNT9��Zj�4�VR�����c`[��!��� 
����P+��Fj�7���,�#5(��%d��c�V��f�<��ȫ{!wsO����G��![���X��ӯk�#0!����7��_Ŭ��84��Q�>r;�V!u��ތM�r�\]�S�7� G��e�m�\�=~��l3Xr�9��8��/-���~X�tU��ƾڙ�\b6�>�S��	��4��Iʹ�))��N���q�������&ؘ�U7'D/C�C�
��h�ܔ��	���;�g���I�T��������������kYk��MR��(�Kf��`��Q��g��y�:�m���D;
@$��B�o��[������^}+:"�;F+�Z�O-�$U(�i1�`*�W	ޤ�(���ʼ��ݜ�8�Y�7����+a	�{BڃW{�g�A�U��a�˥�Xi��JV@����u�h``��
@�)޴�O]]]���	�{0}�#q���yJw�¿y:�rx7���~��/�4r6^]�f-@�d8.��8�e�p���N��L����F�Q������|�t��M���n�"a��U�OFC��2G��5&� OW�E�>2KU���ѓv���k1��ɔ�[�^]�L��&�����2sҶ_^ˇ�Z�ä�D2����D��[5������߳���H�nM�6�1<}��яxA�s߭삥l��������9Ě�$�=bDfx�g��=�.���@�6�h��k3w[��	>��P�l�����Ț ®�Y�q%��r.��}�G������9}Z����dL�/犧�f)�B�k�&������Uu�QR�9'��k�N>(b�ni�����c�V�U瑶`��E��1��Г"��c���Zt��>[۸C�Ѹ8Ѡ�%��NY�ϕ��\�� ���G(��ܬ+�
�8����o!�l"�כ���Q�?%.\�s%���gĐ>^�t�z8�~>ﱮ�٤��3ܮM|�-{�>G�O�c���Pl�����M'�U�g�WbƂ0�QSQ"b�b�f�0WH\*����.�L7AY�o2u�c��u����'-���
����JA�V��<�H�~�Q`m��X!Dl(vZL8Ś�����g�
+��<�豅w�yK˽~g�L��*W��/�Ap���D��e�[^������Sm1��]uj��*u�7�\h+ŋw6�(����*$L�oE]LI��m�Q_;��4	�u�J�00ݤ��x�<h^�c�J�{��Ԑ�����y��n<�jp�_����1�^�5���i��Cc?���B�V@�Vf5�tm�ITPE���b��}cK�u��d()�k y��b>�n�W,^x�1���o���@WDu���sW\���!�@�υF�	�1�����(�X����ԃ�7��(�o^|~�K"�K vt^]߅ф��̋mD�UeX@Dg>���j�Ȗ&��s�؉���|8Y&��5�%��=���>`����h�0��,z|j�����z$8^��LDt׎J�q7&��y&�Gndk_�����hLܛ;��|m�;�NOpԬP;���m��,���
[��m�}��
U���=h���c�@MG&d��P�_G�ه[W;u�B B:|�=����H��j�]jG/D�4�6�~��L'b�&0\�Zl����&�T��t|�פ��w滰[�ߌ,���Ś��~Uh�$K{Thq��B��R|
C���.��h�+P[����sQ�#>���~�e�t$���;e��vV
q�u��[�s�Ƴ:E\�(�����)��_^��:E�/yeX��I��(��Mtڸ6�w������ń|Jʤ��K1o#��^�_Q�����]I�||sJ�����/1�׮(��q^�1մE��OO���3y���[u�&&�-;}��y��tK�`���M���G��4Z+�z���>��ܳ�Y�p]��.�YBF�'�k7a{t=�'Nk:����]X1V������W��ui��|bi
?��y�u฽�&}մ�4f\wR�7��x��3+�3	��ң馽�LY�W+A^?d/E�`�h?(t;�r5`��"Y�'�t�H�y�:���;�ʆ59\�w�S>�ں���D�E�'�����9�3Sf#Ϩp��8�\�N�
�ՈY�3��2���TS�AeuP�=�'����W�zcST~Kʟz�j��b9Qr��	؁�c�m��H$�f���#cHB�S��]zRC���͙�-��dP8��Y�Ǳ?B�,-ŌU��M߭�xS��R?�t�����9<�9�d�N��b� 4�./t5���E���>©߶3:���!�����'%4����?܏��a.�����nЎ����k�ҭ�]��JY���wS����+�� p�z��(~�x~wn��8�z�'9��Nn!@=�KT����$Z��6Lc�o�
;H���qQ
�� �ţ�h��1[mrX��s����}��N/$w� ����:���('�@:"�`���f}�|5h�K���B���u;�U���(�B2�zi�$�{@ā�{S���}���jF��)[�]�n�"z�$WĖ׻�����5���������]2�-/�.lj�T�ʜw�̶M�� ���]a�S)�c��/�)��B!�h
mX���_�8�Ӗ�H�hn[�|\��v��j�_�89�L���64YJ�?v��g��{1�����I7G����H�]���YP]M��J+)��	��Ĭ��*��ϒ&�%��������A5=+d�}葮�J��>�`�=B�c���f�$��eY�{_��j���X!��{��7�v��8��{�{액	��@[>�{35�1���lSh0 �H}�<v�[3�r��{Otl��aOSWU��Q{��h��ZP�Xˑ���C�������B��_*s�x�z�_av���a,��^%4�sN��;���7���5 3�.ĬG�t_�c�w�c&k�x
������
�£��;έ��(�Su< ���!���F!�����̛���'a��F1��Ȉ#���Ο��=n%�9S�3e9V�����t6ֽ)��}�D��5� �'Ħ��)@ה�	��P섹�������^/��Ƥu����|���k��{�r/�|79]�V��d�A-�o�`����x����+����ӫ�4ͽ���k��Dp�sV_AV_��l�z�@�!�{�����b4�[F%�E��u?�$y���	R�R_]����o����Qτ��Cz}�T:��U(�k�5�e_�
J���[u�l��B��$eY�gu�ǜ��Ս��	��\팩�<0\�������8"E�������#��\n[(H&��T�0�B̥[�"�î�n����֍�K�'a�q��� }���e\ۻW������e�ok����߯�9釗�>0#�������I�\�p-��{t�� |�g���F��������)k[�&�/��������Su'�
���A�O1~�"g��j���}��[8W���d�n�U\�I���7�x"�H�9ku�Q�VH�*����׃�]���p�֠�_CS���h&��6�ȟx���k	c
���0��Y	`�a�L��I!\�N��_~#��0����~A��M�H� ��f� ����W�����Biqoq�BѲ��[qwww/�ŋ/���N���aqw׻��?�>��n��$�L����t�s�b2Q�#�X��Qx��k����=y41�%2B����J4�'�C�Q���*�}I��A�LU�0TA-����w��-x(">�ST|Z;�%�u�H+~|�H�V?�R�Xѐ�	����5�P�5��2,JĆ7��:A��1�'�凈[���e� d���F�t.����6�Sc�D����Bwc�@G)��B��
�}����=iKW"�,	��X�q����5�i
���J��Ҡ�Q�,"d�?B?��B�v���~�KA��0#���i�fDb��!LC�v�r)Ɇ����V|�Q�A�c!DB�Iǟ�����I��
���OB��7Y��
b�ؒY��V���-`H2�c"L]j�Яj��$��bd<X�Syl�K3[�C���'md�?�e�u�ewCׂ�9��hN�vfO�mi�)y[ٹ��!����H�j\����&����[�9�p`��c�� �� ��k�����D�C�x�K����T-���4����!>ABCl&Ͱa"@m���5{E<��H���6H�� 2��͝%�Z9�q���X�|��B�5�8]VӗcSF�j|�5(#T��L-;�b	�b0�I[�h��z�.i�c�jw��9���I�Ľ=z�`�E��T�k�����C����3��W�����g�������CA����O�k�l^�.��`�>Wr���`p��y�w�fF(��_ОWH�N�ډ��]�bȅ���G;YD����m����8���V�:Qß��i�-��*�/"�P���@��y����.4&�QwOnI��+y˱�_'=����h�.�K+��>�]�+�$e�(���6�e��ʆM��EЅ��6����D�S'�"�'/�~�^f�	�h�iȤ]�����b����A_��U�H�%��r�׸T���q>�p�=�
���P/��Cg� 1�4�M�
�g0�߿����6�ӿ ��N�{+y�V�4P�R�<�P��5yh����E ���҈z�|1�x������J�{&0�{!��N/��<+S��ID''��t	���-�{�wa�1��յN�(_�C9��!������խ�B�cG/��C"�.">h�X���=a�X�:��?a�D5���&�ˈ�7�{uB�)���b-e�A�.��m`r1�8��f�P�Uw�B7�5��n���M�CY%������2�4r� |�"r�:B ��Vɳ��݃���~�/��9�[�O�d�*��M܌=3�m��ỏ��Ι��aF)�ԫ+���q4�k�b���+N��n��W�ϼ63O�i��Wŭ�Q��M�4;9�
rs:U��jэ<� �_E�3��}��H�ݭ��ن<kk�6A�����r2��D��?I�a��K<�r��2Hl�J]��ʅ����Q-{Bìy��f�*::��6�b�J�G9�b�����؀��U)��:��|�<O�sX�h���ښA� �i��B�6ӵV�v�:���R�D���>�a�:����
u׸&���>�Φ!0��r�� �`�l��`��0˯������2�2���ھ�">'����^]�$�C��>%B�F�Ђ��YxH�Ƽ�b^�[᱋�C�������������:]��q}OB�:00��n���<7�����ׇ�5 Y���9�;/A,��ֶ�B��g�^�Q��`�ػ eZ�����-��e�:�_�[D>g�_�"6
V$r�zy��T�W�R��t�ڼ�HKX\� �R�`˽���8Q�7�/���T���BF0:��{�>I�9�e�%b�K��
]�����ڸ�&)p��D���b����]_�-t����D�x`�;��͢���F�ǚI ׵m} &K�[��z����]��
�Zr����#��J]ս+B�׈���]�_�J&��#�m���n�㥥&�_Z<E)ᇆ�kƼ̩�wJ��(���P�	�E#J�]�l�;��i�@K8�u2����'p8��u}s]`�$ը���p�{j�>�_����T�A�TK���fo+s�'�B�=�E	�;D�Q���9Y"ϒ/�C/1�<�9ĘO��5�}9T�-L�<�u���yg�zRI��r���\���qI(���Lq����	KښF�M�9*f��}.yD>�Y�_f��#օ|��Vq���ej�q����=��F�2i��j�B$2�����8lF��a���9~x���}�w�s�^+��_:�$���T��2�c�/2���,���Q��Ĉ�@�H�b��>>d|}g-��k��?������$���N���dK����e�t��������n�k��F}E�웏ܰ�l4j���D��%��(�ƥϚ��K��H��)rᘠu���`�vz�Kt5ʶ�*F��yDغ���~Iy�x���1�?tq�{19͆;`!$��R��E��!n],��$�}�-&}=�b�J�v��(��r���s�m�|i�wdC��m�o\�WE��l�������ߤ����x�1W��(�z���E%k�����4׋jB9��o�T|��=����#�Rڸ�F���3�txϗ'�.���?(�A���/�b����rMd~y`�da��z*��DZ/n��Lh���4c����J�I<υG���ޢ��)�#4{�S�7��V�۫�N:�k7P��Ø�s.K�v�$i���+����f~��n���m1Czz� ����1�;���w7�E�2 ����fZ��%x=o��z_VhȊ2u!:x��9�뮍��}���3Ѣ�)��ͺ/^:�M��=���5���7���������D��w��y�X������1�iI��� �qPS͆��
�x��T�sM#���$m
�ʦ�)�J�!�T=ʝ��f�9�q�ŋ�Ih��T��b[�}9� �#t��i#3Σ-l-Ʃ�R��c����e~\�9"q��qz� ;\k��D��Y\T����Rb%�W\����i��ܨ��m^~�E;��}��0��Q���Y{x�Ʒ��}�eՂ���b�,#��[L�"�"��2'b����� �M�1g��ݨe��3@��βʿ�L�h�.��ƀ�܁����U���8w��`u7Ԉ$����U�GY()�s�Us���x;���;��0�u��ڼ.QZz��z���c[z0��o���}�����L�m{`,���5��2�ո�򗢸�]�Pic��gr.\�T�����>ܰ�}�O�T��^�Uy���<ĺ��>QI{�QMI�ؖ|BVX��}��
��[P{;�ZW�ɊW�Ǐ��^�ŇT�:��uWo�m�����!x��}Q��fK�?Գ�-�D|��v,��.5ĆQ:n�&٢��h�M� ���w��E��/�w	���4$`KzקYD�d0��;��>rt0�#K���~�"�di%t��������c�A;�[��3q��p ��M�Ǘ���ː����7G߫��dzBK+�eĽE�w[vR^a�tm�LU��1J�ǩ���ma���E�p2&i"Q��u����2�����xj%����t݇ܢ�o�?�&�%pO�g��鿡LA�%b��YеwL-�)DJTG��_�~�E��i"�Ø���t�yO"g�+�A�	Q>ƃ֢e+y��9���uKB�r���
_�������~%;G��|S��V�������uЛ�z"z|�B��x�����t@>�B�rL��?���׽`"�t�E�ה���Y��)��0�D�p�ˏ��R��`j���.{>��~9�م�u3ݹX�B3+�b���� �������߇3Ø*�xw]������oM�@;�Z���1j�ob���Sb!ɨxy8�s>���������˶�v�A;ً"E�wJ3�7GϪ�	���u��j�N�0�ۢF?x=�hD�Y�+#��ޫ�� |4Y'����mL���v�Lo�7Ӓ�1v01w���\� �
z�������b�o�-W
2���J΁�Ԏō!G��=X���BRYC}�`���:�w�D�Pm ӄQ��K���'ڠ�;��I�a�a�|��0!{O���Z��ـ�h�PX�p(��kݠ��"�r>=7�s�+plZ�k���]�ݦ�����)�oUIt�

�b ������mN~����6�C��+�)����5<&�Μ�oGP6�M�6���
<۴�w���n�n8 �NZw��H$Ы��E�I�&.�:��]�<��u~�_�e:��j�5S$�!����Y��1�uwl�����>��'���4:9X�-�a��W�3Os���CW?${4A�X#��A���z���ח�{��������T���/Ws�Zþ���BA��@���U�+ܖ�t��oZ�/�I��5����=���h�k��|�ٟ��q�����,��!M��Ӑd�-�~&֓`�vx�U ������l�S~鳍� ����nu��z�Dzpo����w6k�{3�9b}X��˼�-�^H�����C��+}�&�S�'����A��������ϣ�:<��W�s*L�'d�S���m ���Bk�������;uV|^Ŕ�sv9����7��n��4$��F�i��z	$�:b[@"�p�kt��8�7�ji��l���)R�1�x{ �>>��7ݠ��}�c�`��8z�>��ju�^?�V��T⭅aѧ�ep(�߾�<f�����dԫ6e8(���v�Sx������\�Kw��@F���3Te��i��(QuW�oxL�v	;��o��b�.*���6^8j;�yY���`k��	�Qv�W���(E�oSk��C�y{��l?�ɋ�P�����T��Q�cIVgҭ�����ɩ�������=�X�q��P�O]�I�¡�	��
"f�K�[K9��c�ン�&<D'��?B�=�vl�����)6a�}�h6�|��ǯ'���-,�Us����P2�yG,T�>�U�������+|QKC)�ݕ�����F�Gӆ����̖�W���R�-çu��um�i�'�꾯{�@��ͶU�h[���+��n�AG�;���������$/�)\��T�_A���Q3ѷ><LѥP����r~>��Ir/��ٳ���<zx%���<���r�ɾٚ�q���3�C$y����	�F@ۏv������?��mBy���Q��������9
Y�V6��I���>Gi[�B��a��Ó�*������L]x�
�*Ǔ�{�H�3�N+d��ubX�D��s,���ۢ�%�y�h�2fUC���i�A!.��pz_4�Vb�#������ok����
�8�����b�i�5�>_�szU����G\%?��cK�SV�)�
'd0d����r�#V�ǉ����|^
M�X��_�!&�R��4R�w���.�����>Z�c_鷺i#�@�)4�L����M��!]V�z�b��h3�)3�����v3{CC�vF��V;F=W����A/d�T����罎�4�K�Z2߾�?�y��(��0[���E��ﵙ	��nW�70NR0�W�_��b� �d.3\(�#,�h`������X�"e|�k[2��y��e���Z����kPAI�F�CӀ���)q��՗2I���O��yQ�3j{�ƌ(���%��.E��b�$8���T���X�S�0H�'V��!��2�$<�7y��\��b�u [����E9�P��6Z���c�.�DЏl�>��ў֊{�L��j��ͫ�}y%_X�����7���G� ��a|T�0��,b䜞�z���X�g?N�^њ��D��Z��E�.�Q����a����7[80�^�3m���Q��h�$	t������e9�ǵK�`�A���=�͂���������7���RX��f%p/�i3_�q"?�B���Ma4*�wš���g!�����/Z ��f��|�m�
O���8=�[�W:���]��}S��##gB(�;��[u�(�;�1M�Uy�L���y����+4E��	��en��>8������)P���9�~,���/y�b}<�粶L�e�M�-M��7v������������ˀ+�������T��Ə��n�~w�Q�p��S��T���e���!��k~�˧k��b�mJ"ڑ��;t���N�6�}n�1�;�F��핳�z|f1�����r��v��v��U�1��nN��;�;I���g	Ft��K>�4�wՏ��q��P9�-}oé�!-Zш��qB�y� +�7z�J� ����yMpJ���K.�P�U��~M:+��8.T��E[P��P�y� �\5d1wI�}���%�,���I+��g���㈖�j��Z����Ȥ��7_Yf�Wٗ��f�����o/51�\�����?/s����S�xV<
��J�ӯ���
��%MM�N��oi��h���@���C����&��v~B�>�d�]��J�<KI:���0�bZ�w��	E�9��� ^'�-ɺ�9����������f4�$3Z�_�?I����!�mh��=�c�S����,B����R4X��������m�e�����x��%?Ǟ۷��m�)�����8��?��+��Pes�fV��쐑�JE��"	h�*�~�卶-E�u��Qc�=�%rU���#$��s��uY����~�g�����i���o��]8lπ���KUi=��8\�����еy?f�2ቑ-z�H�bתJo�}{����lzTl.O3Y�Q�>�%��b4�v�8c)B-!�ԌaqKa>�� �ߺ'�
�5m�?���t�Kk*��{�?'g�0��G���O����)_����Q��LN�uz($\��b��]X;����%��:-UG3Kŕ�WdB7��w�O�	��
sF�S3�=oҫ�����5v���t�(T4�M�\gfs[5�Igm��9��a.nm;���*�>j++'�R?e��~��z��OM0�jV�ej��Z�I���O���J��x;w$�؊wW`IbQ���,���D2�S�.�h)�٢����b�H��:ߔ�u�F�ֻ2�mz�۾�q�d�LR̸�QZF��K�ZZ��u�6	�K�MӪN�^�+��A���ޏTIV� b��@��C�t���h:��@ö�����ʓ��@`*��V�:���Hp����!���D��Ŕ�6ɛY�cϼ�x�Y���;*9���2G��_��hq�Y.�ܟ�Hv8<�_��^v��"���Z�e�dOtV�mE�����oR��)�+��x�'��D�-���%K��z��Ֆ��$���ѾfW�$�>��(�*R�RI:���|r��@�ۘ�~��8�"�(Y�l���Yi�C������]�f�ȝ��5Y]ֈD3��w^�!�K&�Q��K��A�Zdr�
���"
��ӎ�;��縥����%T�.6�dt��ґ`5^��H~��f�C���\]��p�2P�;i��e	J�<uZ�5��+3���I�\
�a��QEd$e7���t���D�7��K��|Sz���;�vQR��Y4S(cy%Pt�(}b��
?j�텶�т��^ꔙ֜��D`�j��퉥���,�&N&��F���/4|����S�����Q$�����}��/�q�$14)c�$a��*0'����擒��i�߭�p܊G�߅a�=J9�+b�.�x>Oճi@�CWQ�7���%�a�L�6����{��ͮ���d|��Z����~�N>��}��a�?6��D� ���w��}��dGΫQh�g�(7,�	����f1Kb��y��D_发�SQy7p8��M��J�͸���l�����1�1�&Nܿ�g~\�n #A�R ��̭�U��>
�Xh��l�g�ÃK�W]�_�	=�;�G<�����O���'����b�I��&��$���g	b��XB~ۡs� �Cd�M�eA �E$��/�^&�r�U�&�))	�;�����#��1����o�@�H��Y�{�@��d�)<k�R���_����ن�T���x����~t_5(�'��ըz[��� ����Nֵ:���u~��O=\��n83Q9�e.�ަ5g��ɰ�0γώ�緹	��9ߊ[�pTL�b�Ik�����뭴�N�r�I����毄��A��¨�Bbqҵ������H.��'ǥ�*>w�s VN*'&(��ŵ]q�*�FðE]�=�@s?�Qq{�+��e�;(�L�*���Ez)Ӕh�n�GSn��9�?�l��=u�2k�k)W4a$�;���+���ao�'sr�6�'�������	�[2,T��_�1]}�u�9d���� p1��Ͼ�-�&���w<�I.�w泪�8]y����@�Q�핣˵�#m]ێ�� *f����.#R�z"��z�~#)]s���\��Vi��1�V��_�~϶��;⣓�#�2�����
�����	�^������!scz �%����r��z�!�F��|=�[��yz"��
�["����8*��
�S':�^���\y��~�aM�T���+�;l���:�������%�S ��<B~{���`���Մl1�a�*t����#��1�@UZ�8���Q�K��zimWI��L�S 8���u�1�.��Ngѭ�=o��]D��5�hSz2��[�4�s�{�ٞ⩈'&�;ȗ��h�����������GB����i��؎�s\)fk۱�1�����+�KX�}8�w�y�īw���/��ix��i�T|����fT��J�eR�x5���JA2i����>��`�-8�Y��ĭ�Β�h�F�͍�ƗAA&���VRw�B���g�V�?d�;�\Ќ�8`�DE�n�|d�jZ��=.���-��В9����'���Ysx/9�y��3�+u�gx���h�;��M��kE��'��Պٿlʽh�P+�b���"&el{����vz������=J������<�6Ф�~q��\zr!�"F/	�z�Qf_����C�	1촢Y��t��9�s+Q�<�<�B��_�+�^-_�W<ſn��*�<.��t;���f�`�)vH#7�s+�6O�V_:��k<����rU�3�GYn$̝!6�\|�]�\��GӍꖘ^µD0����Io:d��=��p=ڤU-�,��
�d���r��j�uz>��?���x���3y̡̬1���B��� xӧZ$�{��wqW{�{�}�o��_��8=�k7Ix��9[�&����R�V��J[�Ye�F2Z������!��P�&"�J�UE/�,	H#�L'���*��a-~�UG���?����-Ф���B[�r�}*�^�����aÛ�
���m�uN��܅���lyt�ܦ�ӻ����"���<JA���ҟ�3�=�G��p��I{z�Se!�'�"n�zL��v��4F��<��|�k���c�'�z�'���S�pÓ"���#~��x���C��Iŧ�7��Eg�fb�cj�n~�C@R�t�Ju��E\�^۷#~��Մ~:r�(l/ɜei���	�"��:��w!� 
��#�>�YPQ�>�y/� 6�/���J�KJ�e8�����3�$��B�wE#�d�����X�H�9쓤�W�ǲH[�Gp�pI> i�r����BVS]�i��yLB�&��ʮ�}���
ǚj|<{�����w�P9[	��F����D�g�ZhVQ�]��6Q��f>p'�I����|q�
�U�gά���Q��&Ӡx��"M%�)���4b|~#�a����KKLz��&�o+��\s�'�ZN�q�³ʡ��%2����+�g���=-Շ!Y54.<�JG�4��vzB�����j �
sHGω�l���8�[>_�J�������%c�4狳#ձ�������/�����F��d���7a"z=|I���ɼ�� �&I����9"O�E���fC>�h�1�-���s���4��<4b���<�L �"X��:^>QC@r0�#���Y+�~�LPfA#g��]C>[�×`�_&���,=�_�ꐞ:��}��X���m9XC�&��q�*���{�pD�ô�O���T��ι�V�:�9Q7'4>�$3�T����
%�ٌ�~�.�l��$vSԷM�e��ܳl�8�UC�"W8�t9�����4�ȯ�j�@k�#YD��nj�Q��2ʬ�@�R[%$�����E�_��ݎb;���L�bV�N�с�>7��s��aܯ��ߋ�A
�:�����?#���e���|�;Q5�'����4�{e,[GJ]5�p�\~�p�1�P{�)A_��E�φ�!{�Y�ȧC�*���XS�oIDd�x�J�g��t{v*B$*ltr�˿gd��f�a���R��S�5�I��u�'�%�Z�=���U���`��,p>Cp6�a�|U
*b��>ѹ����g��V�,_v���*/6|�l�׋��B�;0|Z"�2�ّua�tbU_*(g �J4�)K�v��9O��%�aV���m!�*t��N����ɱ���K�l�y��j�.Ǣtb�4^��R��e/鬪ŊO���:���j�v�Nk����]V�)�2�Y?p/`2볬�s��������c�g��oe��'�P<�Vx	a�m�V0s�ʇ�~:8�P��e[!���� /���\�%Z�kU$IO�CC<���5��(�ZC��˘A�GK1��z"���yH�9$5�r}�<l���{�?��0�M#@ՊV��Hia��0��$P� �b��Z��E�A+%���r��i\�7�|�s'8pȋ�A"w�b ��K�5�`p�[�k��W>���%Wu�(�С7U���I��l�%	0�������[ߧÁ$̝�ja}�m;�9(��@�4ӂ����=�_�B$������kQ�Y�e��E����M�9O�!�U�F�wD*�o�!�%���X��J�/MfĜ�HxS�=����T�QI�L�:��N�U26ӄ�r�D!�z�ؿ!nP/�7BQ ��Mͣ#��I���кwm�<<��U��`���I1y���m37?��&A���oૻ�V�����7�Μ�HA��� 
"ReP)�D�6����|��-�i��Um�$��|��ql��L2n�?��޲��.p�9H����[R����ԷJ�(b�tL�tD�R|;�=��QlX:Qe�g��^���C�����I�V���L�o�8��n����L�cA�-�`�fAK Uq��Uh�i�~�PI���k���ߪ V
�g.9��br�����[x�\��T����+d���6�9�f�M��`C��{�I��5�[�1�l0����(Y�$�� �[�\=�r�~��v"��xq5��Ⱦa���@� I�#�wK�D�y��P�DA�pA�Cء�Ǥ$�o�W�o�&��������K�W4�`('���«������
7�~��-)��������lEE�J���/�9i�N���II9J��Q(�F���"�9J6�oj�I�ʥ�~�
�b�G��J���v(��X} !jC���r� "}t �I8�<p�'����ua��=�F�CL
��O��J�f�uST\�Ҕ:��PHS8D���q����5��?�E�!ʙ����h���~�_B9�>@�����
�MNo�-�b���?L�@���Ax�
�u`K���d���A�0B����Q������8a���Bd������j������+��Tb�H �{ߜ�1ě� ��&��}�,���?6��~̡ˆ2}	��`N)�	B��}t\��s��M��nZR'SF�TiH/��O����D%�)�ӱ�e�6dҁ�:����@��Br.J �q��_��!7Q}0�5\��!(�-a��7L�<ԭ�ä>�/�ǤnZ���G >�<�Y{���� �Y��5?,JZ�*_C�x�&1��j��=�������+5_�
pѴ�y��n*<����$�^z�33ޔ���B����V@'��`0-ܩ��vL�(w�N�~�
WI�Ac�9����P�D���6BV@�����XD�37$�I������i�4M`���pe�����>����tN
D��{� |�����.��͍�n���`m��B�
W��ED'��'�P@���yz�2�2ƀ�����0y���v�`��I\LG��W��H�_���8/���(��#��B+R;����o�s�V#&�?�ג���V#��X���='ix����	~�c�m�L�܎�mz���B��tc�`��#����x=:���ٲ�c'�<�{���~�!�\.���H�+�{��^��ݓ��A�7�۬�'FJ�Ӈj������{�F�.�����Q2e¯vwnI��WT3������є�1�<[��M'� ��;(7Ǧ�t�B�.[��GW��g윀�Tңʩ�]Ym4r.�G�_�yj���z�y~[L!�r�̄1+d��c�I97���54�@�m�͓�l���j|շ|��|�����3p�b���Fda��\�E�m�_;+|F�9�o�qj�7n��O*���C�x��'=6��,�;4�/Ag	h8e|��T�d�.��~�Q����
��&~����|V�c/�1���#To�(�\	Q��J^4�z�W�Orҷ/-��3��c�[� ��4�q����v<��^5�1�U�AH{�g�ڑSVV��n�{]eu6��D2�#^�%�usQ��'��#���Se#���GK����ƈ�P�2J���a��5V�\�Lf�g(����٭Qx��b�Ƚk�9�]@�V����I��ĳ!8=�;���}��6t�׭���P�KV�=�ي�;���!-D������"���a��o���v㸼��ݏ�{00|�FN�^vU�YU�-�hq�BΜ��=��{:v���dH��i����VSu��?�-�x�E�w��}�OJME�?���IE"�g��=�Rs��s�4c�����K�q�TtyѼ'Z͏:�n���ǟ�������xp}��KDU,<梉''���KN� $�M��ښ���a�a`F�q|��}���^��[G��~ȳc�7��އ���6���.�o�s����ӿ�$�j���X�`���F�n��%ב�	儆�6t��zܳ��?�o��ħ���������WǗh�y�bb�*���.X&��>CM$*@�\|����K!�IQkG!B�B�+l��!��o���jыa��Q�s �pV�7
��z������_A55�3�R ��&��y�Q�х�a�G�I�=�,�V�͍�`]�!C����u�6#tҷK}��ϯ.a�'W�wo���l嶩��p��
a_��\B�o�Z��[C��\uCfIJ�a���������o�P������~���I8n�%uc���ip�i�ӈE�^�z����Q�~Q"�G��&���XxH��O<>튟o�u�V�c��m����2\l;����ﶅ]b?��e��C��=�4�$y��L8D&svɏ�$�y\�b��E�9 ��Zot]7J:�T���c�yI�>�_ut�R4�p������ڀ=no���p3��
���XM�ODC ��p\��"�K[ё�f���d8�4��	mI��3���3,�Z��h�ր��znM,t�|{��Z~FQ$H����D��X�yB~���9�f�8�Y�x������.aT�ƥw��p�yR�Ǻ��Ǽ��dE��k�2��r�F�i?�k��z��1�_"#N���H�~5�cY<�.�%Ňà�����àOq���o�n�;���Q��[��5�Pѯ��\ҵ�Gk4�z٭Y��F����$�j� ���������'�"�����R?����o�sA����I��<�w���4�����x[�q[�cO7o�-�[/M��§z]���b]��N�୆�Z�����B�ʺ^��W���,g����o�{^7������^mz�/�Y��|�w
QJs�N(+�*����i�{�y�~[�����D�*ʵi��Y�D�*����m@.�4�=7l�r���~��(o+s�M���a�b|a�RVشq��_�~/�������g*Z���B��\�I&���!W,w�w��Ѱc�2W����Y���@�;	C�K�����-"���|������z?��ꭓ��)ۘ�2���s�/�쀛�	��ڑ��Fà�5�T���2�&�hb����߃��t�n� �>x�'4��\���O�(-�S�pm�QD �-�J�L�\�����'+��7i����׈t�����$U�9\\Ӹ�V�,��i��?��/���BI��EO�4��?d���U�V@:ã~#(��ƨ-Nz�V0��X������Z[�����b���#�Rb���t<4"�$�C�yՋ�\�R�9[�嘵,)��i(�m@#S���5��)^OiR@{l�̯s�|{&����M`�r'S��1&m��3;�����(���-�lY^��p�Ś)?щ�Y<��bS�T0����=�R��������yEr/r���?���JBԴ��R��}�n��ʫl,8$X���Y,ɡ�r+��cf��`[��&�Pt�&ǳ�ƫw�w�Ik�K�r���5j��$�pG��0�_6�ڜ����(i����8�����' ҹ�z�7^�>�[���������#�vj��^���ر��)��Z|��
X�! ���p IaV�N�w�<:P2�������(۔>�����y-�!/{N��Hd���k��º��E%4A+�25<�����qg.ԃ#V���Տm1ufs�.L�	u� Iz4��
K6�?;�Z�C���|���|[�~�U��6�C��m�7�֞��'�C���E�(y�����뾜��|��!�Kh��'mj�9v"��b��\!׼��ǀ�T�����N�.<4���>ed.�:Ԣk>v~>�Q֨8�/3/$�c`�tϣ���,��
���d���"��Z^�f�@`sl i~M��fC�&�8�c�C����ilS��\��gxlL�_��{Rڙc���� ��)�C�ű����=��򼀻:���0��kR��q�46�in&ѵ���*�t�4*�:�ѦjC0*�A��ܮF+�+}�T�˛gXd�*JN�L�� S9� :�W�v��%^y:��K�
��8!;��`�,���>���Zu[� �����W@�pP"��0�7�X��2���n�||E�B�1�K)[Q���ȧ���rK�!�9�l��r�I.����+N���YJ��Um_pf�T��u�N���饮P��a���/�n�\��8��Y��0������[��=9; .zX��Mbo?���׻�l��^�Hs�9ģ���J���_ΜpφegL�
�x��<-��=.�1N�M�5[Ɨ�e��6־@��9�Rg���?xT������VӬ3��0H@�Ƃ$�;��ƫ-��"��0��d$��C��r��1�g[��r&Z[��k���}�`�)�>��ͅ�k�p⎋o�T$��m�u�e�h5^�/���>1i+�+<�ʧ�W;��f)�d��:���2bC�=�ֻ��@�CĽ����G"�ns��G�s���,��q��n�����s�^�"R�����~ᒨc�������V�G��4\�Ҩ_��c�kI��U}n� �_�7��]l�s�ܾ6a�q��C]r4ۣ=���3��VEE�e�%�kF�	>
�I ����-sS�W9��`�
�z`k�C^�}�r�L�2Rf�M��z��_,�k!���we��'�C��xk�0�!L�ˏ�/��W���--w&O���b�uǵ��""8���q2�$�6x|�i}n�
������yI=���.���R����*�z��u>���ʎW�V�pެ/�."�t�L�h��X�9�*w��Ba[���i��O��WXG=�q��7y��<q�J��~�a{/Q��b���rc�39��4>C��xw�y�Ų�<27^p��+�}�if�;�!i�|�����d������ ��G�"G�Q&������4�ޞ�75�Jv|��{Y��&���l�kq)��9>!�ty4-��aa� b��͛��YF5˺���*-��V����/����x�/x�ʏ3[0޿�.�Bӽ��Ʃ4�ч5K����WǺ�#������t��i#.4ϖ{/��՟t
{����|�2p�8�H4�Q/�It�f8��	�Y+�^���K�"��om�*u%f;՗��|��
�<*��l4�2�3���.��r�Y��f������QT��:2L&�X5�`"O>g;h��m��xZ#:���;�i���̋�K5_�z��y=�U����:+�pഭ�	>4����@O��0���5�E&o��a��0�Y�p*������I��������:h8緬���yFwI��G���K��|\�?�0�<.��TK��D�D�6�gK�H�H���&�����^�x|K���>��&��)���G�Ti�rD�z'�=�!,L�7y�Q�	L��h����LU~V��=1�o��x�Si�N�y�j��h���p,*���>�kw$:#Վ��E��	��(l#w�Em$^ÅZ�T����8�i����ѺKr�3$n�Z����9:��mgb۶��F�4N�6�����vҠQ۶���|o�������s����s�ٗl������E�d��'��5�J����q �ܢ`�Z"��`?�@�`�/^���=/��i2y��j��Ʃ�Ν|�:?�>�}]$#:���Ƨ�Bc<O�o�*ѿs�����q6a�ʎ5��&�T ��(�O�Ypnh�,`}'�ݗ�|c����z�5Z�tO���
Del65����kf�?���V����iڷ;@�����p�^	n1�z���_�.�����s]�f+�Y��

7�Z�y�gÆw��v�/�f���W&��߲���f����on�L+%~�F��q���{v���܁��V��7d�
9Or�����=��b҉"y	�[%ϐI.��0�.T"���3��ǵ�kq��S��D���Ӯ<[0-`18������Fr��8!R��̋��Z:����M�I��A��z �ѫ
��������۔W�Fx (��~�
��������nm�(�e�	:ʠ�ј�F�/U7jm�'m,DV�T����X��W0��Ƌ���
_U�"�e�1�|R�A���lM������H����1��pl�y;���z�4�+C�ϻn�q�����@������<�h��4��qK��'���:���[{�;;� �X���
��[�����_�r�"��,��D��w^����f�8[Z�I1�e�c؟+�V�įM�e�Q��.XF��y��n+���`�d��
��.�)��v��>�KX��|�˷[D���%�9$�h�B�ɍ�"�,�
��`ɏ	^��͞-�m ��F;thk�����`����m���A��V�P��d���x�וx�C���^mv���Q1,wP������{�&Sɚg��#v'�aC��%�A�JY��)��]lWU[�Ů��@�w�s�+kx����?��/A���PD5s��[S��n�A�`���P:P��F5|������K�*M_]'R�Q���Q�!����:�^�b����.����`�,gl�rkn� o���!�7I�O���
u�-[8=?�o�4�����NE���o~�E�>�z�i@Z���ٝ�Ƿ�Lհ�5[c|l������ �o���YK�K�c@<����V�"b4'ðS\��_�A��?dY���-,ث����7��m!�޻"�Q�s8a3Jifi�M���A���l.X��u=9I���o�?��r��}�/� *F�������w��x��_�N�O��F3?��'�U����%X���)�%,�+M�O��P֮�|%a�����!������%%?P�9�e���@�<�~�b��q?�����d�����Q�f@ ��\��ɉ[P�ʩ�3�kf}Q|���a��#�f�j�uu,t���b��O��K)� I���֙ыx�f`*��m`�q��=��aX�˳
����H���`�Eew������+sP�MW���7j_ʗ\%.BuZ��s6������u2���G��%
���߷�ѬIDv�Ȟn(6>�U�< ����B%����Lr ����w���4��E�W�Ĩ�t��,Ѷ��iѣ&.�q��&#=�0b|5d�C���v�6��M��!��d=���4RH*\}>Q��U�3"As��2��/(��y$5�����g�2��ն>5��M���_]�����|���N�2�Ot~D'��ڮ}�<=�{��g��\�
�G&�1�`_'��J�ZW�阹N�xF���	�[Vc{�ً���h�r�cv�n;���L-5�~GrĖR/&�����:�t��X��wqC�F����x���/����~|�Uq�!&�7\��$R!#2Y(�F��lV����}Lkj�����9���7Ԟ�:�D��ǳ1��J8Ǘf�������#Mڅ��R��y����=�0��P�!�p���JZn~�$����9�J�Q��������H�k5�;`%
uOxNT��ɔV^9��͑���������Z�q��pޞ���.{oO�Oݒ�~9:/<Ȼ�e�!��:�����p�y��й��Bmm�;�IB��\8�wa��x�����z��#8ӆ��*�Ŏʊ�Q�pfS�V���k���*��4c���?�O�U���p�>lHu�8ӌ'A�c�)s��+�1�� 9,��r�z�OZQ@X.	�ZO�YUK�n���6Z^�W�jh�m�|%�O�|?`���mf�<+���(�>U ��\������5�#����#�	(jHk�:�������G�11���X�ϥ�IY�bj��_d٦VKO^���ԃ_�m���V���5�O�R��T�q��޿K���70�;��Ǔ��dQF �*�&q��ˌUo/1�/�	^�W��6��6���f{�z`e�솚�B�w�S�ԏ#U�؀��O��f"\1s�}�m��B��\)�s	f%9������*"�nn�P����ד��]h«�c;nEx���x�Z(/���e:��_�gHr Bh�A8-�i��f����H�i�?x�� t_AL��Qh�R�m�����;�9.�y�?6a�WVV/2�'''	�4��9�p����N�D2i�aN6]�e�A�e��@u���зn��S":��;��J��_t�$�9ƻ��Y�b�"V�o��Ytq�����J��G"����ӵ/$������}�w6�$�۲�`��,`��y����C�Mi�6 ����#�X���J�:����LN	�m��"�'>�٪������`��-+��)9��@r��--����"�!BJ�oװ���{�M���ƿ*e��'q3�o�Tɔ�_j��DH������QSV����	�HEhT`}]�q%0�p��,ezD#U��N:�3,.�0ګ� &���X?�d��=	2��F���:a�aEC^�M�,�Baw,�yoG��
C���+5�b���^^T��]`�>���1�l^"��:�#���烞L���O�aaaMVУ1��; ���Ы������U��+�*���m�J�b����ۛ���v���B��7��M'/��a�ނˏoj�$�EP����X�<��?3/~�i��x�*e'�hA���7>��;ɘ�/ �>*�v�Q@kͅ��"���T�����2"4N�D�!.g[���Y\D�	�\PJ�>z8K�:��1�m��1��19jU$"�FK�I]oJW�尿�B�}���QȆ(��@��w�vQ���n�V���pp:�0-Ӽ�P�\�I�˱�9|��5(�>Mz=n7[8ڮ�ɢU�>TB��Zh>�Ǒx���n"U����T����pg��ʧ!��es���Al��{kSX�����m��>5
.�oo�5:�\���*�;C)���FU�2���F��N4�4�_�*�ݮ�P�w ���Ꮣ��ü�4NF�����Ӻ<�/�,����-�<M���-Ւ����h�?��c!�Eؿ����A��]��7.r�f���sE��cge�l��LݫXӀ6ն�������^c�x><T�w��۾ͲD�ײ�J��ƖϬ4�`3(L�Z6�$��i��q+��("cNur4�r��s����	C/��u��W����g7���wa�m���}�e��d7��nV�)�H��;��$7���U��r�&��(B��*�VݎBs�"��Gq�Q��5>B�@�)R�i<��O�8�zPE�z�N��z��RJ���o����:��7���o�[GR�J�a�//!W��<�|Ɉ�[F=�v���`��y���Ո�K���T��>�A����σ)�_s5����T�~�#��Z1��C�c#����m0��8���s�ʔ6�"#Zg:�x'I�N��G�X%wiݯa�/`KK�F��Ր�Pn33�i���'7�\�O�%�}����m�ߺ#c�w��LoW�+uD���TO|�����1�!�C^����]�|q�$y�2�R�)�!b�)ck�ρ���l�@ӀdV����"�ݨOb�Q�T������!.���6�F�	�:��" Vq1���w#rG\�D�RFe<)C1���=<�+(�O��Yހ���b(3���tv}�W��nLG��Z�D��$n���G7��~�Ъ��Wad(�'N���U�N�q���[��$�w�q�K�O�4 7n9E6���RD�礲)�T����o]��I82on�i��������uw��ܾ���#{���(�������=k+D'�MXkDC��AAA*P���D�R����$��c��Y�o�$=�����Q<��𞊻V%��x���oN/���o�7�s�rЉ6��Ӆ�=�����|�7�AZ��q}�)]`� ��J��+��a�]E6��$
��ll~�9P=�w�&�B{�c�A%/� I��Y�9���M*�}����R@�.�
њ���>�^�Ϣ����M�'\�e�f�k��ߧ:ςF�Ń����$����6�{��xe9\��(W�9u�q�?1��������
�h�{��H8k�ө�����=E*�_m�g��	@��=[м��B$��e��^8'������`u�(���o�	4ayktM��ͥ�c���u�#d]���.]�u�������o��D4�0�	��Ƴ,ړ:�j��w�ȋ���[���My+9s�.6Í��>8鉟(`�z���N�.t�4���~��5�#u�\,���&�9 ˷7�������;�?O�$:7�6�K&��Q��ahc�j��@�d����YO[a+��EsO�ڞL���$t��,!�Q��?���
�q+T;�k�����7�r�,��
|��`��\0 ��5�<ܱGq,g�}ܕ�!Xi<5��o��������9������ڱ�hoˣ7S�_�㓍, &5jcE&Kaiྼ|���{�Xt9���}������9C�踩���Z*��	�N䬇���Q��>�"��B��޷���z�PjT"����ۉP4��~��Mx��}��#�[�B���#��l������ ��"�YǩD��wǣs�����=�ڄ�k���v��0@�(�zi�＝��qڜ���}ܬ|2�~�\��^�_ә��䌇�@ ��t�5�47t��ȞL
c"�����N/�K���3S���O#Kq��	�2�,����V�8/�/n1�7�&(H�T1���\�r�v���)Q�,�M�9�\�0k�ߊ2m���͘,�o�Q�Kd�� �l(�w_�1 ����о ��,���u��K9K�u����4��M�jv�����ͼ���t�E1K�-��2��-�G��\�˄��/-��Fŧ����$\�x�C{뮱��h!�]X�y�,��Ɉ�?�)�j_�D�c.O�LM6R�|��sՠA����@���ߛ�3�
4�y���H�ʄ�7[1~���o���"&n,ǡǳ�2��.��3�ۛ�O���Ԉ��A����!k:�VC�ۄ�2�gqJ�՞d�b�x�X tM�
� � .݀hy�='C�m{�z�2�ĸ�.bNc�� �P�ǳ���E�I���6��]��[Nq0J�$�՜L���i:-��	Z���7Yt�_�L�7��[��
Xq�k�WQZ��>S�2ReYBׯy$C%�3�'r�Aђ�^N����4T:��G ��H��I�qF5��&z�3���۫���4Q}7�I'��X�����yǒS-ܻ�SD���
����>�gC�ٞI2��~$���e |�[>g�O� ?'�b�j�A@�YY>a�k�
2������E �.�����N4j~L)	�S*�k���x�?��NY��|�g�=�b��٘
zb�4({���у���S�ǐ�#�-e鏳7LQv|�kX�FW""�j7j~�H�[�V�_��#�*�
�/ƴ'.Z:"��"��;�K1oUh����P��z����H��,Tm3�xX<�񔓫g}'i�:�#� �} vp��Ԩ.M���b��4�D�r��I��!�C�!���Ք��l�I�`$����JЅ�c�$�;���w�t=!�&](]����pk�O2��]�|�UR����>㔻ݛ�e��^Pq��V�#ş1~���ׯ?�2`��N�m���u��D�2��+�3-&%���PH�3�B!���:���$�����:�B�J=�s;jCk�b;�
��nu��3�J"Qe�F��%ŷm+��Y��%e5��Ȗ�dqj>k	r�B�vtl��g>I�i&v?��x�#�-�ŸH��j�R��[���A���u�Z���y�D��1rD�%4\�������Z���s%i�A�D���������"���BЩ÷�#8bADDTI�Dp�u

2��f�X����r�'	)�h@����&N��,����a�!GBah�3q_�|	<X�����T���m� ������^���[��z��
A�HGBI@�d�E�`�Gh�7X9<�\��@|U�=�$���8�[�cp�-�L�������cȏ$�)��?��c(�B�x1p�X>M"���d�`�w@��[2��,��S@�~..�0�1n0�� f#0A���v	�""�8`�s ��<�`�	@� )	oEZ��,�X��L���/!��Y�"v�G� 3a��9��� ��g(�A����$	?�&F�@$Wq��NC:�'.ů����(d��E�M�E�I���W&� ���ǎ�AQ�MC�95[�"m�}`@sڠ�9���ϗέ� �Ɨyv��|^��6s1��R� ?F�>�Z�<��lE}�o���������u�$��T�{> ���((BGk���=��q��)(&U�3�ܕ����W�j��p�Ȓ��P�BF����`T�� ��B*,=w�\w��W���t_�����T@|���Z��+(�s�̧����oK�"7R��A���������j>!�C�|�Ə;P�˻�Ԕ"�����t��p�R�� wU�?B4�8�-"u��� ����P~5���u�V�_R��Zi� q��]�'�z����Õ9{�!�������跶*�	�\lEo\�T���R��-����xV KU9Yy݈�cNp�w93������M1�s��V�Zk����j�[>8B"@��nNoh��9�9"��SJ�..��FڔW$Т ��䳜~R�ѢE��.�4��X4Jn��kw�3j��Q��_�����.���Ln����D]�9�Y�|X��kۿ�S�W o��nȀǃ��o�*�	��A#uӱ�m��{Cm�}'*U,D}���6����!��_!J��G�;�~�?���o�
���o>k�4��|r�����y�JӹkS�����C�\Xa	;`+ŷ�{,���?+v/�ꝟ��CFzn��%�
]�����&��]�H0W���~[�?��@��v��B���8���t��%ra�ƛl��N��јϩ+6ӊ�q����TP<���g"��Ôb�
���g��U"z��#�d��cv�$����E�����s#���~ˣ]���e��*Z�
�v�)��v�LQ6\1���z���(��	N�M.	��W7�vO�l���sFª��m�\��3��2��vD���R��	�1Cw�G���!��S���F�qf�u��Ҟc7��7�=>I�R�����;1Ϫ���s��F�#Ud��0ѥ��Sl_�zY�ͩ�����a��ӳ����"�/��S��݄�u��d�F�b���g������!����R30�,�JD�Ѫ&AqK7���� Z��z�Ă�V��fi)+#��:I�7d� �R�/��7 ����8�Wq�������nӞ�ܤtc��v��9GA�]�'��'N��������y�އ(E�غ�2�-�Ղ�����(`��G_�̌O}��=Kx4��d3rF��j�Q/��H��}���|^�̻[�`�T[a�f���r+!��F��a4�d��M)��|Dzmf"�*1�f�'��b�?�{�+v�x��j
p�h�D���G+��WǕ0�n=m?~=���J��b���ή!��h����z%����<|�l�_Y^$􎠼A�c��e����-��p֝����=���K�et�)�n�|u�k���Z�s!i����.�ѕ �p�W1�!xzb��C�=U�@AM��Y/��7 �-3b�o�M�D��8�n�%���ΊJ@�kf��� (�|�+-���(^�:�S7�zq7g�^��������'������ߎ����Y� Z�E*����j�����qz�|���Q��9f�ah(�����}C�5�u���d�=�_|]J�,�@pFZ�v�*�����F�(ٮ%e���S������K�ۮ���,����Dڈ{�{K>-
�,��
�;��ƍ�7}ܪ�+�d���!�"�X��X�����]��j�m諛>�*���kE���	̻���<h��~)�|M'z��>�<����x1�[f,{i��=�rГz��\�����Խu�����6��>C����t��f⪮;�-9�u{&�B���)ku�đ�4W*�=���I�h��j(�~zֵB;H�M���c���}���PQ1f��
�M,�-�Y&a1�(s�zO�z7%�ћ���Wu1{`Ӌ�×*V�v���ʍ�g�_ȔN<~�؝J���{)��ߙ�����Ek1%�'2��b�tE�~9�O,է��Y�~�vU=���h����[0¯��z�#{:��Q!۬>�&�_Ӟ_P�E!W<1L��ō��1~����̻��e�y�Ux�.�.��?P��x�"rϨ��me��Y��-��,#���й�2�z�5z)���z�6E�#��%mN�V�p�[�r{36���,��|��<�C�bPV���vs�������v?�I7�W9�k���%qX���O%�Mò�8&�fY���Oö�����6�߿B�x��B��0��gv�2$3��8�������8��7�.�)�(\g�BF��$G�e6o��۞��^�k-Z��5ý��%ݓ�"�'Q\�(Դ�q�v�M�*��(�\�Tx{U�e٨RFZ}�И"�hi��[?��B�����t��h�����B�q4�X��x�8"]j��6����<��?�a���>N�W 1rm҉j�.��0��#%s2�j�n�(��d1��b�9zD��l��:�n���c�1�������t������N齫{�yLݷˠ㊧�g�܎>k=��v�Ş17�(g�I��ê�v6wv����Gȶ���� �T�n8�+Vl�+���t��-�T���i�N>��?���]Z�*B8���m�ⅿ�ZϪ0����H�=�k���һ���l`�r��g��t����`��I��fA�VX����-�(o��r�c�dOl�#��dϛsU���
��^�����=��7�����z��֊vI�&�'��\
�Zm�i�K����)U�s�d��f�>&��3H�BL�)�A��ܐ��N�5h�▽�r��r��(�V,�v�]P�~k���w��� ���}!M �k����㛩�)ׂ耡Tc� [Ϝ���$uo?�&C��Ӄ��kv�¥�pX��ԉ*��j|]�QZPbJv�8�ZvQ��{��k9DG	K�L�t��˓�����E��.����	���P?%�2��4-�K4rQԪw�2��R�~�e��|�.��3|�2��뜫&�)X��M"D����rt-������e=-������?��>�	q�y�K�Ŵ�o��鸖3p&�/Ӥ/��\���I�i_�7D��d��ׄ�h�u�
��Jp�ĵ�N�N�� |���R�k��S�4\[-_&�U��pJ��������{$�O�~��AG,$)�Jܺ���4�F؉�U4E���L��Xby�V��������".aeʣ�P�ᚙO�=��=�0�?7���{2�?$�$�1uͼ%�=p�"i_���,/�V|Ye���d�FLw`�c�\ҶS����WR�K�XX�|�˪�S�r�r�`���;Ү���dX��Ln<[���XmnmՉ@_����a�:��!�}�ٽ��(<ff�*�g+�xo�,��K���ٱ�#�J��`�_l¨+����l��ڢ�
R���-�)A��LZʑ@��3u��N@��\LL^f&b���LP�~���Pt<����ߑ����������\���iG@3�QFz���_���(����EI(�U��j"��\�eˊ$�Rlw^V&c�VԖm]��6��/��<<^��M�n����U�1��%�����m���F^6nɘ�y�|��~�;BAE�f��3���[k�C�w������4��)6I@�1�筡FVy 7;��[N�"�7.�.-� �1���a99�CF�2/�KGJm�KU�j��m��9��h�ː�%{��Q�mO�\f/����]Yclȵ�5`�Nb��v:���ul?�����4u��pTK�KRaJ�:sF ����$̏�l�^���[{��6����5���[0�%ڿ��6gR�oo����{(���ܖ}�[���R7��y�Л��4Z���Ǭ�~@�����}�d���7�)W�n�`��C��6Ӕi�y��u2b��H��(�1�	1.o��Q#	=P�,�E$�B/-QJԥ�*s��d��:?-sEr	/u���ڢ��w(z�qAYB%f���v�;���q���0�����7Y���3I��e킢D�����U7�`G�]��)2��j�{�W��/��P�`ꔲ�n�a�M:I��JH��-n�:4�������}�H���ܭ(��i�x�H����^+�݅>%�3�E;�k�&�|P�l��~�܎� )��M�������JWŉq�"�e[���{�v�����a`�� [Q�tģ(]�G��FB\��$��@v�ue_�
��$o���EQ�ǜiv	�eZA5'�Fw��~R������\���e-l,��
���}-���:��d�JXD'�<4�
�?_h{fO�U�Aź%��6PU��'�O0$դ��_+�'|�HJ�ms!�W4��C{X�<��wb��rͫz��O�|�A�fv�A� ����=;�ߋ��rͲ������rhfD������x�Ҍ�[7�vQ�7�`?�'(2o?KW�8�Re͓G�D˘�f"$D�&��tbE(¾R?�^C��m��v:�q��Ī����ϯ�ܗ���p��)�t�J��{�R�d�Pb��$�-�T9��kyP^7xKW Hu������ ���>�.m�>�hf(fI-�)RT�)&uj�{}1�w���4C�B�#8l�u8��;�E�Tg�+D�\(N�Y(c�^��98sd�d�����ȡ�@E�+@GdڗBsa���X�5dH�&��>���������i��$"RC�7Эڎ_�,�h&����+^4�1S�F�Aa�h
�7P^�2������0l����7c���D@(�]+��qC�P����������$Jo�$Ni��5*�ɣ�tb�8�T���~��4��j�EoĬ-q��r:��6ndE�E*(�J���\���������q�:�8ј���բ��b�8tAZ>�����~ևH�������ZKn�O=�l���Ox�Y��Q�4F��Z���e��Eڄ���^FA�ݽK�1m��u��m�x������������w؃F���;T(U�b���`jb��9b�*�ub���[k��*zDJ����L&�3����7�W����U#'�Ǔ�l�m8�9����)�*���3����*�k��}"�	tֺ+I)��p<�i����]گ��)׼?�#J��/�Ď� �i���g�k� �Ӌ�v��`�cC!Ɩ\�eO��Us#��ΝQL,�\��Q��1U��n�nYz�x�&SV���ߵ�{@S �~~JN{k|���9��?S�Bp���]�M"�5���zRv�:U<'��r���j�F|��܍f��P��}�Sgn*R�~��N ��[�V����mH�R�`ݽ�@��x0f&|B�W��Mo��H�J��B	�����%�*�����}�;��R�+��#��)�j��H���2l��+K�S�ٔ�������.�f���ȹƘ�	��W�%�H>l�\���kq�Z�gȨ����e�X��z�t�����_v��|�{*jC�� �,�ߍjfC5��a��:j���y!�*�bbU1���Sk!Q�-������ƴ�hɩN�fS����@XNċ�`�ô�XDt!�J��(%�4G���ZGo}�,v��I<�Q�uaz@鐔��2��;f��ӛ���N�:�8Iz�Z�"�mGW'�(�r5Hr�lV
4 �բ�%N4bA���#���?��IB&�6H��X���n��wy���î� ����$!G_��}Y`�(���"z<̒����P���[W�m�ۋ�1}"8��q���@9�S�%�	�&B��SN�l��i�-�Y"��D6̱������ɻ���_�n�?`4���P����Sέ���C��K�a���](�v�R�		�E��V�_�*CG��юֱ��|�Y=�(a�����E�6�y�8$����l�5���2�HtLKvQpZz0{��d#n���h\�Q�̓[Q���2{0�����ɲl�@=��` ��dԶzS@%�P�A���D�!i=H5>����A<8���*C�mx2��Dє�D����+Њ��(��;�x6J�܋�.)|!Z��?�G��p/@Z��bL� A�K��	�	:�|\(`$���u��fL_d��X	1'&TJ"�)P9Ef�\d��t����y���ʻs������k�s��b��đ+n��rB�58��GS���b��L�^�.TIzĭ�fi+��$$~�nB������2O������n��en8N��).�cf�J)�W��{Y�}��x�d�5�(�"SZh������5G}8�~7�\~�	^�`W�)�����O+���C�Ӯ���{
q�ڠ�ωF�:"�N>��a�R�+�R��ն�����L/^+�!�Z�~�
�I����D����¦�f���~�k�K�{=;�`cz����e���
��U!&�*�`��}<�c����W�0D<y�3�X*@���z'hyBBf�� 3����ࠇ���:|�օ�.��K��e1��
����}Cn�#6�^Cr.PE��)!�D̯q����G}��Zg�����<�w*�����t����Y_�R9ݺ	ǜ�}FN�3��ǚ#�?�א�><��N����9�cy ���I�'�01��(����g�w[;���S����aJ���g��=�O絮�L[3;֜��^QB̬�1-�̭3A��XF�dE�;�Ui]�g����:u������Ev�+�zI��Z�JM�R��FZي&]�<̞���FI�&����ǟؑ�ڠ��1v,&�@��4��ȾT�x�)SF�:Y[%⠇ml��\���]��H�3�2�G�%��\Y�:0��L��N8���m���3K�j�}��Yc`���̞�+j��֙/��E��H�Ӽ��0g�=U�c;cM����NE�MF�����G6@�-NFF����/�����g�*ӡ#^�RN��Kl��DEE!���Zߖ�|���	�ֲծ��,	gJ2���ɏ)�L�U\ω�jq>�]��!;�3Qo𸲭���VѺy;c{��=4镻��T���>��߾���x$��Lr�,St (��|�O0�Ɲ.�S*�'�gi�~|@���*�}m��V�|^]V�Em��������v������cGE[�<V;X�Ukj�6"Ù��߿�JLR;�y��^�1��C��kGOh��L�Z$Z�M)�ϓ	��)�&Eү_ݷeS�ݭɋ_�,�s*H���Z����C���2��mN�hP@g��AX�a��X�����je�3侒!ݙ�R.\ޠe�@��ɺ�Ao�f�D��p�L�`e�>uN$�a���p�'��#O_*��V;�~�Lc��GP���m�;��$���8d>�FT�����$�0?H�����|%Ĳ����B������%�k�?�E]�2;R�W=�C�9ԡ�`
1[6�'n����﵍@��v��8r'��%M�g�'~�u���W,���-FQʢ���ıy&|޿lR@����~����Je��w/�}������4�I 	=�R�l�/��|Q��w�[^b�����||�V���UM�@ڶFT����7Uc�i��W�O!�(�޼�S���'�����7�s��f,���b��U��GuE��޸��	������_T�8�	ь_�y��_S���Lq�"�G��h�4Κ�®��!��*�؁�z1f?�(Х����������+ �:G�������㙶8U{y�ਔ͈C~��%��O���h�����ւ�/� s���5Afe�B�J���M��l��@�������'-(�PZ6�� �yOOc����/%iC�ү9춧�.ؐG��̨��`�M>��_^�6��%�3�q]�;�3\���6��d���~�#V���Ћymh��6K#q�����C��Í!$�?u���"5~��Rm�G�k�m��'t��zJ)HN�HW{<�u�Ax=G'�ʇ|�}tt�\�􋒲���NU�bПN�K ~��g��)L���I�˫0�i�ˁxG�R�܊gϾI��}D�F��aK`����=�0g�U���f�2�)&~��c�IԻD�'��|ֈ��Uoo~7���c ����(�/d��H���6+1��^U�@F4���/d*X5�d<M����Xm��dbn�)��TY�s�r���8ؘ���i��L��X��x|(�uj��g���v�q�WYܗ��-1ډY�D�}�1)j`�L�}q|�VO+���wX�k���#�s�N��&�Z�o�^�ĥ_I�� ��w���y@Ũ.�]Cs�:���a���T�g6��ps�|2��c���	��7��L�5VH�E�1E���~���D3��4���`/K�7��#�T��H*u��n8Wm�~��SQi�_6�_{z�j�7X���RiĿ�9.=rM,̭��\�Ǒ]�f\�(t'R��ė���P���V"�����Zz��T��N�2� ������7�e���wbV�@�_��0|��e}a��oVs���ܓILoYa��7�f��&y�W��L�|,�E1t :�k��i�CD��Y4t����"�\�$����<T������9��:�d�uM�L��ZF��R�Q�l!݀����P�?���N�}�0��L;��=0tL\!��^I��'��(���<%2��V�t,�h�B��Mt@���$�|gý_P�*�>S�{�"�x�߬��QT�V=sTK-ê"{�16IG*%��;ʞ�R�����ݹw��<_w��=����c|B)j�0�X���A�3���"k�s��Ѥf$[�c\zrso�[�F�rXy
����"�����x��.�������h����O.!n�����'喭��-E��K��8�<��̱N{0�ge��<S1ϭI,iB����BOt?���.Dwt��+���|�{'��_iؔ�w�����Mga*
V�\59����"n���3k����)�#}H�{h�h^ۄEr��< �n(b��{L�{zDz��j)d׋����mVqo�/-$n����}��D[I>*���2e>@p;���@�7�؆�'�H����g*��t
S���i��f�Aڽ���� �?g����_䝽�E<�hO�IۑؓM�V��d��lK���b0�a�_�bF�W�`�Ա2}����ej1@[���X`�B�¹
g��==q(�)"���I�{�r5貞�4vp���s��h�W_>V��ڷ�����hؚ�����MBD���{�1��y��O��U|�]���	c#٧�8��Cp�dC�E����Rve3���ձ�r�5�4n蘭���?���#-2�w�z�祣��i���P���բx���p�Z�}�t)��(>���'Anǆ� ��"��o0n�L�g�dr�R��b�$fн�$_���N��(	�S���5glc�^/az]*+�z���҂�k���	/[��cPC#�2)�Ԛjv�YXy�mC���ʛ�����������PG`v��AM�$��qar��d����h���ؖ��5QiLZ=�Tn��L��K�#(�ǣ���:g�� &�B�rx|���V�=�}��*��i�7v�����`o�t�ì�%&�j�
mu�x�<�M,�)�QhR(��p����[g*.�j���M�m5|1�A��Q?�����y�ޱ���c#�;TJ}U1�O����]��#��eI"5�%�}��:��:�Ӝ2u�����q�R�">)x�҉�9�����s��a���7`eI5:�88�+Tz�v.b1.�Rk��)}�ݧ^Z1`�����.��Y�n��3�8I��e�� �]`�N⍂\�	=����m��#��%k����y�;o���q�?L%g�EYik3�׆\dk(E�H�:w&��$o���C���u.N����:�E/�M,89��u:���K���m'�����h�9&M����2*j�د�����Y����	�&kd%pC6����]_q�"|�'��A��1we{�
�_�+"�������1�^��6��؊�,�W|.j����;�g�t]��;�m��c۶ӱm۶m���8w����>���h�k��uUͪ�Uc�0f�j�Գ�++��¦������|�B�0��1����Qx5����{�RV%�-�컜.�m��I�PL���ga���?v�b�8�jE괈����v�2ҙ�̻�����l���N��������Z��4s�#�~+eU�f����H(UK�5�U���u>��Yr̈Q�����R�$�`�ik������6��v����T���|���bQ'����i:0	���f�7��Y���Kic�-iW���Z(������g�J�6���e#7���c�Ob]- ʔ�N���2�兛�f�j;3�*�`�d��d�]���b/P��BH�:�qo�O��2���w��[1ܺ9ӊ�9v؝{���^r��4��x�oBš>��A�%YX�ϕ��uTu���M��O�f�6��,��'��/*J���'� ?ENt�
.`�[1�N�_\En#~�$���t���s�q�E�g-�Օx�� �7ѫTt��|I�R�u��DG-�s�<Tr��vue�x��69�#J�6�+��n����	0}���@�德!�>�E~/����A�M��.�\�*>(pm��8����Y���GC����U���+��rii_MЎGx�꤈��Pȝ���6��%D�����O�'��MY�G��������lT���6�/�����J:έ��*8o%@`y�6����5��U�QʢQ��;���v�]�6��� �m'y�,�Fmt�D�{�y��)R��CDYH�m��DAD���HG��C�Zrel�&^Eq�������nY�z�|����Z����a��WK
�d%ɏ��2/��H���Hȼ��
���(ִ�DGt\T�H���ge�@���,��o��0WM|�q>�y�D45��H��)���I���zrR��&Rj�ABيI���ӂ�H�+�Αą�_7|�x���e�e��o#UZ���EY���֢�U�w��i��J�z�,Lc�B'a��ݩ�j���꽗&xj:�3&Ԣ��=����E��"��Ɇ�����.�u�j��[�1����>�c��?K�ψ�_�rt!U�7ߵ�V�����?d�$e6D�����[C�.�6%�A��I[�v�zA�N�r�Sy�����5|�������J��Q}��&���(g��<����
��j{d�U��J���Fk�Z��ݗ��{uh.��e����N���վ:��|F�h4�R@�X1c�i	|����A�j*�@f�����w!KzUx�
��燽6WsD�ۓ��j�@�^G�A��sX�4�ox���1�{?=���݆LG^��Й�4H??�^I�T/����2��Ad�1�%�/�p�e��[�����"�]�Ґ�ز�h�<涷/���y���$#�h�x�3�_F�hѦ��}4�wha]�a9�bxI;����q�D�,�c��}��=/P}. �Ӎ�q��p��Y�l�������=��T�S��������gS�/�n��
�P���~�����N(<"k�����Zɔ�	06VC���V����K%�򻴲|�z��C�^���*�K�e�g5�����o���y�L�����'8���a�搑 ~h�	_�CN�(�ص��� ɸ��)�U$���?�	#����e�I���p��P�E�
-���Y�t�W*u[]o���-ng�u`����%�����=����cF$l0�&v&�3u;=��GȋeG��5�򈗺��n�ԕ����"�L�T�Mq`�^��iZ�j���"�+���p�T�k)	���Rz	��g�o'���_~"���;�@Ȑ��k�F�ЧŜ
�,ҍ�L/x��h!�@�D��⤫�!�@!d��B\���AQ1q43)86�mi�.��
�:v�7���r��*Vg�T��_M�@��gV��z����ە�o�b�S�l������ k�g�KAڒO�;�jyY��)�x���{��A�p�T�ϯ��J�Q����[��J!d;~>L|[c*eG�<��#4� �(#��U!���x��W��j��j,R��罃ꥅ�'���`�+�Đ+,�{W6���G#7���_'����L!�GH���$
nA����"�}+u���~|����q������|'�IXz�y,FrC�e>E��P�G!���'�k>Ɛ�gʸ�NR6A����ϰ��`�W���4%�����3g����#����06/���@���.y2�؄�$�M�x�L2�?��2�&�$�Z�\�S���&�5i�&�Zc�U��`{Y%�!PN��PSl{Y�6K���!1��/S3|�����P����
�����I���G��0nTW�_��Z-t6ꐈ�=.�{[U��V��P���4w�1��5EÑy��Q*0�Cicҫ�v�����a�X���N� ~Ia�G�K�tx���٢,�Va�%���i���0���Ős�!��N���J�ZQ��Q�e\*o�9�)u��p�'��J��T� ��ɤI��jѱ��(���a�a�������!�~�tLA6*���ݚM�h\�,g��ߔƙ���2�ϑhV��g*��:V��"�K`����V�X~+���:;���M����:]��<�-U�q<O����hw����/
���%��o��(%�WKv���4Wtjy��ر�|죻8�E;v��
��)L��.����_�_��~![c!�̄�#[���7�K�.�RE&	�CHƔ`[H�.�L�O��L��Ib��(I��!��/~^c�asl�6G��f�v�z>�|ݪ3)����}�"A7��S�����mU�Z�Ҙ.�@c�1���%�|��q��f�MU#��a"��ӣ\�6t����X��3��~�cS��E@�X���+�PG7W�x�`��͕n��#�ۣ��7p��PP�tb�ʍ�s�}���tb��"���a]h̕�%���;�&�nl�}]���dc�^�wPI^`���X(k����^�e� ��*�l�����E �8�K���{�Z��ȅ���@u\�T�g�.Q9k�L���Ӫ�+ěԀ�y�����~Lb�$e]��@��+t̃\��Ĉ����u�Ɓ��J�@��"j���p��d���F���l9yA8��a��D�G�Gk��ʒ��z�>�ؔ��9�C��~���{���n�d����(��6�t����o�uQe��:���Ľ��h��	��1�%o��J=
F�|���cǯ$ζ����S�ϼm��梕1�I-?�n
����?���u��Y~��rm��������h
W�%^k�v�'f�M�ɀ��;��6�z��ᒭ�AC����J��������(z��}�O��F��f��.�e�=2R�Z2��yT�d���"��)��x[��ǯxGр����ج�\���`6�� j�f�΀KF;;)�/FlV{��M�zHt%�ź�e>�:Ē�1||�ٌ��E {�.[w�����[%��RR�2�^S�P��Qzj�rߑ��Ġ|9$�:|��r�A	7�8\���	�r��.��d��^���}����w�줖O¿������b��/� ��p��z��\qYD�o-Q��78��,��Ǫϐ�)�D]� �gWݾl�@tܤ����z]�#[����� ���s���t�:2�2X0�Ov����� �k�mn^�y��g1��@�Á10�8�`��oMw˯/�;�hʡ��d��g�B�&]àQ�V:�YO��u��^��֏{{�OoA���y�A�]ة-p(Ao�瓞��j�V����m�(�]��0�<NJz~#������J��;^������G�`W2�8��OCV�L� �q"���Rn���@���$��;y:)��c<c��f��b��@�)-�v��.ޡ�{R#��iC%�����BY���T�����3<�~��(bX?����8E�^�lw�����-��@$?K���������v��u/���F�� �g�.�<R�av�j�������'KG5`P]ؖ'ʭC� �]�ͥ�G�[�v�{G�/M�6�`EC����As���Qܓ�������e�'��_%���`�KZj`O�Z3Ĕ�l&ŧK�U`+h2�-��}����u��e��e)f��k��(Wc!��O�10�q��u�<����eνm��I	iz�ɺ��{��s����J��P���#�wldS�^���#Z~����f��N���$��F��ZǕ���Ĩ�2�Lі��.<Ώ��|X$���EϢ��_3V�VI���Rp�*��A�v�����3���|�L��Z�ϥ�A9W�ҟ�l�������~���?H
59��;����7��	1��ll*4"��:0y�0�M��K�b{&t�H��V^��3@���wr%�v)93��E��p@���BO�K��?�:<2������7�P>�|o{~;پ_uB�U�;ݚ�����3�0)w`���:U�1�(�n&U]�̞�{�֡��
_�O�_al���XN����bA��k�8��L,I��/'��c�gK�ƽ���q��G�ķ��ȱ�BP�ڋ�������S��^�;"s��*�f�jf~��v>��j����p��QQ"+v��c0�3;�2���ñ�hI��&4L���&JaM�X�
A`.:_*�6��$'+�k�?�n+�5�:F%j~�'�R���b �A��!�3�F�Lk>L<)׆�u�T=�UEɎA��lF^N992�u�ߦh'Ɇ=��P����&rUN�{^�b���Ĩ��B���������"�6��x�l����� �|��������z.�����Z~��B"'�P��<��,�H��O�1Gg3.N�j�����xA��L��Js��y� RIP7�X4߅�0{ҙ�ԗ�YE�&4�˯��e}��x��i�C�P�o2ؤ�&�&�"\�����+�A��^�>�').���L�����9���+�C.971�N+�yP���Pr�j�ڒ��K/DxCG¯_��a�Bm�9*�ܧ�|�$���'����u���Bx��x�x��&T;^�����z\��
J`m�H���x[��$��//~چ��B��A�<qM�����a��zV�Ǫ��y�,�PAE�*f��í���mK�{��\��	D�hVvW��l�M,�ʱ$Eؿ*ks|t�$k�����L*�Cyi�5⮈#&
L�Nj��$ɰ8N�$K��4��q%�c����`ol�Z�t�dU��&�^�UT�>~KU��x����WΛ6�]��l�#�h�g�q�&>�1Z����X1��F���D�1�e���K/�^Z�3r?ÉD��t���8�+��%TK��_�%�i]��1D����B�G����~^Õnk���/�u8d����ƙ^�,�]��O��4܆�ZP.��� �}Y��c�9՘aLbka���=���=��H���Sq��\)�,Us\j����j�hҢ�ST������Z~����v�O�9J��������0آ����N�I��3���?V�tMJ.Wn�rE���p��)-O���}ا�9��R*B5�%hdiPt��*�(d�]��d���\g*����^ޯWL��z �ﺱXcE/c��M1cs�y��7�z�9�x�[�߅$�J��?�e����[�:�n��g�
ozzs��{���+��]%E��yN���)�	�8~�^-���A)Ɖ���V��P���z�9�IF�S1�O����&�]���c����gTd:�#>w��e�?,#��(��"LM�3R���O�����x�O�v`E"Q�u��BPp]��RN�_�&CJ���� ����Pf��C��`�{<NIe[�=S�5E0;�C��!K=ET���[^��'�z��J�dNyv}�Ev*��Q�F�b�}9�x����y���^)��$��j�8K�!'u}9�lB��o����@��S1��z��x4��:*˜�bp�`�c��H!릵V#"�����8�/2�s�%�ʦ��jp%`�#/���"���͢�������҂N�X J��W��;xJ#���0�T�\>{|�L�?r~�nr�LE�)��JN����A%(�˩���IKu���`����fN�lq���P�BO,sC������h�6�)��%uO���O��g9 ��
���9R�!���Y������E\�w��I8�4d�l-�wp���
�Pk֝��_�"��&D3����w��d7��Ta8s�χ	����>���9J�#�É(x�E��aD[�̖�H�[cH����B�����y��T�iI.�ă��ײU��O�f�(�v\��aR	xeVV*���.Mנ8�?����b�'H��%{�fo5V�
qE�N=,
UP�����rY]1CC>��CO(�VS�S��������V�D�W�'�M}�W�{�t�Q�@��O>��Ԧ����� mMU�uڭcX�
3��
OW�8��9�&O�%,0\E��?��@��8��~v9f�~B'u�SOf�����έ����I��8b������IB$[:)�Ɛ���^U?��}#�����efxi�;	'[�eӰ|�y�&�@��&g�]�m��Y� O�!y\��N���^&��˵�t��cEȎ)S��˾��CUJ^���`����ۛ$v��ApJ"G&�W���O�p)�O��Z��4��2����TU�o�����w
��1�Yq�(M��H��o��I,�7>�w7��A�������Xb��d��kH��s�}����$�Dۋ�����_�(ƿ��h�}���R�?\�_f��bzM&��,4��y����T���8�ا���H�����,G�XO�f7c�`�����on��%\��w4(Iٜ��&!�}��W��1�9���>*��z���'�(���3|a�:y��E,���R�G�d֣�,4�j��߽�W�yS��B�#�m��^��^vwۚqb��(�M=7�Zip90s��4���!��#�C���a�L��lo�sK3@/�θ�=30�ɭ~�+�����ӄF,)-�J��]�6�<�5�����$57���!��c��?���FaK,�P\ԛ���ꓩ�6!���m���;�NtnZ
;nѸɆŷO�m[fn-�$�x�c�8�)ت��˭_�o��B�4��a���]��QO$���@�:�i��!?�wP(��'M˔|?����@�K8PЅ+{TH��
��~�VU��j�9sY����O {dJ禾J�@�$��K%J����v.�����گ���v���������c4��d�� f��i:߀dz�i�u��}�+��2����Sy���-f�t(�����\鍰XpvC���|�W���[��z��,��_?;�;����h��h?�9J�L��71��i�e��i�?���[	O<>�.����)&�G?=������Z*�B�\ɰ��㌅�Z�ie��V��(cn���s>P`I����=��CHX�>���_Ic|��ܥ�H����;��7�J�(t;e^�\Ni�j�.9"?fHe��=�|oa�7�$ؿ�t������X�����������.�a��0�+��Ҷ��E��;�?0�N�����N�xHKBh����_%I���2��C62��1������͋qETI����"��Bt����!#A&h��]�+�x��*���#��~�;�,�8�	S�X�^l��N��!�?�M�@�V8�MySS0��VoesV6��Z
7��|�8?�Wt��#���H��շ�f�db.P��T�nsȏ�3A/<g���ʇ Z0u�s���Rdu�{��i	DS	�Q���S�>�z��|z���Qo�S��4Y��-��D��erǮ�>�{Le�>�}�Q�R�P�>R��&	���v�I<�o.���1L����~Wy��s.Z`�Z�
z�����
��5d���n-�}�-|E�j!(�nD!DC���H�!�)�*�jPS�)�O���"�|ຟ����[9�tv���:�.Yk_���D&R��m�ȉB�B���Cr`�]��t�ᾰ�_�	�Í��gWk:T�(���8�
��F[I]�f7���d�o�R�$Ŗ��Eau�c0m}�Y��7ٴRP�W��Y����o#�w�+M8��$��<��@:{N�`�å�KXI�81Qw��6��-�P4�WcfF�j|�]����&;��s��j��N�u��7!Mn���@f���{��Q���(����7�W�7w�N��`Ö�jڣ����:�v��n�G�:������U��`/���.D�Y���H�ۣ�^=�_�`b����PҰ��j��5��{�e>�e	@ l�}�A�q��g��]�褧�@ݥ:ڋ�O��(7(�P�%���D��x��d{�M,t���T�FP3ڛ
�4SzE�2��Iw�#���X[�D.ӳt��GG&4T�ϔG/f|H������������M�����	-G��c;�͝�^s�>M��KQ�9C�#0�gF4*����^�E(/�E8�Y)�JJyVf�4[����'���sI@�U��p�=eL��t��Tz�z����U�!K�Ňi8�T��׵hc�Y�Ӕ��[����UQ̲�0o�����HE��i}�s_B�� h��G���-�'�����"a���"�uy���J:�8�~���oql��m�~т����^��)q1���+^�����YjWV�7r�JK����ؿǕJ�J���L�j���a��;,Xگ+� `"�}u��7�}��!Vs�秉h�O���O橩����&��Ҡv�Gw�׵�Gr,Je���3� ��K���N�F�_��P�����[��n��u�8"��1��
� ��0�P��S��ZAb�+p"�@��ϖ�>�R=�I�E�&��ԭ���dw]~[��[v@���ވ&3�AS*�Q �`��l���.40b?a(����x�G0a�ްd];��<L�	>�-.W�Ls@��_�����B���B\���9�8#�M�8��R@�]�<�cM�$�H�N���lkL_�x\m��>4�9?��ωk(%-�ND]+���uz���'�<�i�����Y�D����Ւ?-T�4��fNO>��*K�N�9W���UE_ޣl�0�N~�U]�P g���e|6=Td༷�=����^�����RA�@��Gt���*�����ݾ�/�f�E�a̫ k0I�����xh2X�r]��o��Y����0�4Q��Vt����AP�_7Q�Î�or(�*�zr0L�|�"58y|��\�k� 83q�g�D2M�w�!�ڪeR�]
�!\;i����U��.ے�O�LC�n�J�A@��D�U%̯٥���Q�a���E���K�$*�}��nPlk���2l�g2�Ûd
����ϔC.�b��T������h�wT@j�7���5>V�ĩM�D.�f�|�u�.�C�3P��$�q"~���[?����ר�2�4>�:vP��IcX�`1�ӏ�����ײ#�
�u@��1H�p�T�������ٓY��ߞ��}��n"��X[9��PU/zo[����G ��XE*�R�7�������QvsY��k󧜈&�\��g�p���j,y��Rq��jЅ���\ǎ��l�?<rGc����-@��éj�(�<�I�k�h��c��|az��q���m����Ғ|�ŧ���Hl-�5I��>z�	���*�^ef����6½���;��R�2�_�����ͷt؄m,���/�UMi���4�͖	;��6�'A>w�y�?^-p�EA�p��o�nE!��>�8c��u�}�����M��*�||���o�1��#�5&P�4���ڑ�,&,�G�0ƾ��mK�!���Z�����w�AIɉRy�9c׵]:�Ƴv9�%�в�>5�Q@��5(��'�[45	��R�KHՋr wޅ��w�:GL�B<�b
~s��=���˂�jB6�a�i}E�:�cH��]	k����?��VL�&��[6�"��H^J�C%�@,�q����kb�9�M#�����6	�^�D�z�+�Z!�4�I�~�Mu�k�Zx��..��GE���W沧wx'+��\9��-Q)�\�������)�ȂE�҂�Ѵ�fu\<>��^0��ww�!%Kŉ~�UI_��e��aRSN��b�k�*'gbk[��$I+�~Nh�ڋ�B<�6a
���`	'��I�.���A����b��Xj8:���٬��sj�kuS�o���]�c^�V
g9[�s���b�Fނ�	�Z��O`��]�ΠE�)�P�U~������	4��8/EI?���|\\\<�DEE��pчh@��V�*붏����Hj��ш+
�k�_�,bHn�7���w���܅Hh(:�y����2D��]���#ό@QK��a�)�|b+���K|Q9��7��o�r�o$£��ap~�(�_��߇)�kh�`P����n����D�J������r:#���-��b�KgHR��˷�XK�<�%��M9������7A"��o��te�g<����	�GֲR�X�޳k�2G���l�K�j������)~�I+Ot4w�ÉT4����r�D�BV��o��IN�6���_�l�ʆ�y99ق*�#�v���r >�L���SrT��\uQ%6�Fޤ,��� ,d�[�`a�+��s��A�Gq��5�R�f��X�&�{<����y�$�X��{�D��.��r�#�f���V�S?��ɶ1'<ߏ�9�� @�����XX��\�/ %�C�8x2�qݜ�#�TSW0!��QgD�)�}��w�(�װ�qB��g����r�t�%C����Ln���{H��ыR�b/#b��stŎ]�^�54�P��/X�TR�Cj��$�����Ȱ&�'q�S9*��"�R�d��|��N���$/(�>�	h�4Cܘ`WQ�Y�=�63��{3ĸ�� ����=	�����V�urFc��M���2! �5�G�Qά�v(��Fc�;I���wsty��E�������J��B �5StQM�N#���\�v�O���"+������^&��v�ʊ]�_{ns6�[t:�;��U��52Ƽ�I�;$�ƅ���Ky����?9-S�k"A`��X���O����:Y��I�ȳ�G(���/2�t}tەΒ�q�� F� <Mb�W�it������f�:������Z�g@������������oh.z���@�?��|�x[�8*T�Y��ެj�ykƨX�L%�F'��Ea��&[O{|nq��S����t��1�����Qg/�-e܈B�[� ��'W6-*�M�(Q�'���[2���X/s�a�
�d��H;�KX�v��K`�[�U��a"ݖ�꧱4gh(�;k�4�a��=C�@-Hb}6�=����f=2IT��� tPK�ż�9z1H��R@��Rt~��ٍ�����I���>`g���t��k�@#2_ZFzW�k/�S���`���0�/2�����]���ͦO�t�cp�:�vGa
�2'KL���]��@=!��4��� �D[��J����d�W���k2�c��Z�.�.�w���x?c�FP���c��=uݚ�@ ���	/���z�=����RL�c�`�\ZlB`�$�����#���4v�av� ��4���F� �U�2����~*��߬�qw
��S��������G�G˺�[C�
I������Ե��e#G�j�B��4�Biy? J���쪓j������3��i1��pK��(ҋ�o�lA���TG+wʢ�-[�D��ް���,���]s4�>Z�D� ��j#릊���P�c�v����d�JU�a�:���� �6[��"��bs�UPu���׾q��|����1�41޷��#Vƨ��L��M�N�.��L�A{�ƴ'�������2m�z����Sn���m^UV��.	ZrI�#����)���p�tn��O?{X���_�{�x�&�Y�pߧ�xn��h*�2EJ��!W�.�ϧ��;`���������6ӵ�4�o����C�Q�Qi����[w�GN�"�J�oPX�n��<R�ЮM=o!��wɀZ����>M�(VN���J����4�5�K��;�4�cP���\ A aЄ�ŃϞ�d]&�/�{ϩ�����n�&S�t�fHs@���ء����B�a�3��ӜT3�Vx�:	Fk:"3�������=]���bM��xw��;����ț%����"�b�>�p=D����{��Q����{T�ѐ��?�f�	w�??ZgHqv8s��9_}F8�6�Q�jO�;~�F�:j���j��s� ��joΟLc%����כ|"u����2l�[5R�!C4(ĥ{o| A�1����?�f�5FhS��IEC�Q��k��DBy|��2�LBC�6�£fv|�pЬ��ʰ́�7u�@����f����� �^�Ƚ��LK�D��5�B"=�h�����}o�n���Q�
 �i�����&R�#ѫ��S o&��q��.N��w���F� ��&׭�=d��I�drd)���(�g�r��:z�Y������I4��!# �䲃���P���_�x��[���e
k����A�X\§�h"�������U�Ǐa)���Hg�D��K7^�]2K���)(Jm��AF�
��G?���ұ�6����K>��e�j�R�����}Nqg۵P!����x�j�dXCb�E��N�}��%>���*���RU(\�O5�����h�O]`�
���2�
�06��{����f�]7�Z�I�$����g7/��I%����>ٽn?_�I��+�mo�����vb�ߎc6�߿��P�w������Ei[z�L����w���%�F�wYU�x��@�=X�L;�E�V�Ɯ� � ĕ��2wP���V�(^^@�.s�<�n�Zy'�sխ]
���c,@o2�����]��
ԯ��=�!�4�šX��R��Y�sօ�MJ���#OGFiԉ�"��dҖA<5k����nn�d�A��;��ܢ����7�����vA.�#�Z�)��DmĎ��j���51y{��j�B�)���_đpG��:I
�KhW#0Ó]��D"������)A�0h2T�@�TA��)��5X)�Kh�ھ��Y���PeZ~�IּKu�7�pQ<�N0r�L��а��@մ���5.�Wr��>	�|쒐�1~�R�NO��S�I�����8�P&_�7�T�r�H�"�P�OUr����M���j9�	ݮ�f�a�w��dBM�k��^BVXR��]��|$=��=��C2�ޔq�fF�G��Ѕ�(Na���Ll��"�H֚��!����
Qg?Z_�-I��dn����`��+���	�{A^f�D+�(o���ټ�!Y�O�%E,��@;�<���$�׊6Á�|M�wvކ��HJ���]���K���c�$��p��oc
}?�BChш���#����������1�����q�
Z�4[�
M�A/Ys(哋��\��]^p$����L�_��yC2q��P�8$��f����C 'g5��@�|����w}��A!Di�x��8�&j,��5�D�λ ᳧�7R�J>D����&���7qQQ��F͑7Wh�Um�Q���5K�̮�i-V��]�K���K`�8S1)^~����]yD�γfn��hA}PCT�l�����1����L��۩�o������ֵ�3�ի���s���_	�{���]�?G�sB���O���➽e��ѤÁB��wJ����8�G�3_�_F7����p��&�`&��5F�K���ɧ���,����9b����4���T���m�V��-`��7��:Z��P���-�ž��A��O�K�3��e��}Aso^��bh"aM��ғK{"o�J��H''!r�8����7`�I4C٣�m��?@��no���Dy�q�.1�>���d�:k��U.���6�����9  +
f:�~Jwo��1	��A$ΰK�Ե���D:Ju]l��4�P&�����L�5�L.T`laZ6�֌�)��r�"e�}�*��]��J��eP���G�d����H8#�0l"��b�v�&��6�6��Q~�E��"be_Q�=$6��ܫߍ�X�����⪬��b��������]H����Uc���f0(;��r�=�[���=i|�1��`۠������)5	����MAn�$
�X^V�v{sƼ�Z����$�Vߺ�Ic,�49d�hnNFECS�x �ə+$�(}���>���r��e���v����+�WX�L��VTSh�{G�o�!p�N`��V*-�ƺ�D�Ba�tP�{{�d{��+*�����Lo$t� q��t�3[�uZ$��e�)ʼ�}3����%$�5%½�p�P����~�q�檵�i5?(��z�id#"�r��$G�Jz[�U�Y�ǾQWO��]E�f���_�g�f�\������P_�4Y�Ȝ�m���#���,��z��ӂ���"�%%!A�B�����2��V���������C��Q�Zz��$�r�"�vC�ᐔ���Wt�eѢ���H���K����U���ʔH/�7Ȗ6�Q�v@%~X�7�!�x���ȅ��^+�^��������e B"����)t��UdQ�� $H�7���q�M�4�!��r�Dv���yM�&fO��N��&=%Y)��A5�����mO����VQP���U
Z�d�*2�P����]N�} ����{Z����׃ך���1�7�b�J|����^U�c�;.R�1(�`��3m��V@��GM0��4z)�ӒV�~��:��.iʫ��	#���W'��ʑ�!w8����}{����y������/�K]%�a��bZV	J��$�0�+w�ˊ���uN�w����t��L��i��J�#hq�m.��\E�s5%�`����� ��0pd4P�z1���π���؃��4���]�x���d֞���E=;	}S��g;�/�1R��珘���Av;��|}f�$�B�شT��m��@�t�r�-Ї2�6%g[���H9t�h1ѱG s�r��\¹����m#��m;��RaSs���!�x��hz���=��s�=)�u7����(D�]F��1�h��C'O�T��[l�V��`"�7�&�B��v�.��	E�YE��oy����x[hVe�B)g�6�%��w1�Xwb2�R��B�`��8�ͼ��T��MP�*Br��V5�)�"�3�d�dg�'��'c�B�0�����<�&6/[=�a��!���R���.m���g�vIvm�}Zw�ˊ�I�T�8�T
o�Wp:��Fq�5i�<������x<=*��t`%mkBo]&��3X]Ƃf�s�:�p�?Mt����L�pTh��ɋ��`ϼ����|fb��_��:�"u]�M��Fa@�� ��q:�;o����?q��B=qW�B|��b��ra[�����R��0Jy�u��6��nۮt35��n��Fnzk7���0�l�]���9�� ����n��ImVi�#�[M�(�M�������( 7/qp%�����s��	�#�H}�w�{����EL�e9��+�9�����H���y�k�u��ohhe����:'���̖6�U�۠�aIw�o�n��!1�E�5��}��/]׬���U+�h�6�:���N��1a��Ր{]�4�z��^gtֵ��ژHII�<:�a�<7*�(,�����t�.9ْtd�74gЅ�Pw�ߓڡ��WԠRX�r�
��=$K�Ms��s�t�_'�8���(�b
)���^�Z��+1g(��4��?0�`'�V�.�'�'C�ߕ�^\������zp�d�9�׏A���=�/vK}8��?���8����U���m����P.
�(��s�|25l�{����K�|��t���i��u%�@C"����!��}�O(�-@���fS��k9Λҁ���X���(�les����7ps%�qDa����T�n5����q-��o�x˲�Zh�]cwp�Ԙ/!�!_��ŀ��3��du,e˭͠�ʽ�Y���坙��A|�Q��������"��u�ydK����Ds�����6�9��k^��0���v\�X���f ��iUte8p���]��,���P��	WjȎ����'�hm�?`D�w!��W+X�3-�?�-:�
�NFW�d韉�+>���<�xd��P�ː��v�XF����5^x�Q`��H]m��������v��B^V!�5��AH)ޛ��<X�Z�h-�ۅ﭅�W��?ܽeW]�-
!�����[����8��%�;wk���w<���q�?��j�ڵkW�%s.�����,����Z4�����V�ˏd����,�_���0,=���J��`��wn`��r��t�.+s�\�����l��E��ɓGj�T��� ����]�[�GN����U}���Zv����sZ�೰|���_\��{4@ &���_Ϋ���wQ6���"�_ңa��	�2�-�#&�r�ݡ�n�ȳi�Ưa�w쉭�ᅖ�pTuwu�i��1g�b�X3�h|Q Kq'����������`Ă���f_��{S�%�z��R�n�D*�Z'�O����O�J��`Ƀ}���_��>��vS�W֋�ǀ�t��KJ��i>�����G�P6�)�B�1`1�R�kQ4�����@�gno���|��n�㍯d5��<�Kǥ�5g6��Z����*BMģC��umɍ��'�K��);+�����W�  8�&�+�7sr��tE)&�m5tLۧ�{1���uYq�t+ҽm�����FKZ�)5T"9Y��,��*d�U�Z>L<������ɔ�9�ی�nlr�?,�ۀ�9ؚ��Z$���RL%8�=����/_9��40�DFrl��ܟ	�2[,�����"0n��'b�z|��^R�ϧG�f�eF�����S����x�՜�	雱���t^^/>��O��]��{��|~��w��3Q�ӳO~g�wB�Kӎ�uĲ��w��N�����'4\O�3ն)3R��ꍮ�x��Ԍ�_�?ʐ��)�i=�Ln2.݈����
o��i'L�S51��\�#�9�ĵ�Uv0���
#��ha\�y�}?2�u�^-ɔ�p�˱ɪ�Di��-qn��Q���7#g�n%���
'��;����`��M-8\=��#��]�T�kqi�Wg~�,���.

E����;��)/�u/!��,Q�I�P�OQA��,�_Z�Y�AM�H y��KQة��T�<��{�8��k%,��U�ғ�I���c��b�O�Q��+��2�Qo6�lP�y���B��+�t�y�������_��y��ϼ�Xۛ)��M ��a��.߂�RC�rWڱ��@č؟Q�N.�R�G�g5�;��d��O�x��4LEd5��g�>Z�J�jGJ8c�C��Y��%x�;��8���h���=�ϳ��\��bl��ܻ�G��k0�,��_7E=@���m/��6�kӣZ.y��@��j��g`�	�����D���;�\Xw�H�_	M��E�L��qg�o8��>}��>�r�(L.(:���F��M��h��F�&��]����R�,��A,�܃���m���;��gx�>#*jl-M+����"����Zr��i���C(��@����� ��h�xX�o<+^�><�7�~����Ա�Z��3Q7�'�Hq�Xtr�-�#��D֍ z�����I�D;��,�&��K�o��9��6#�m�)$�Mk@�ӝ�k"���ǔ6�So6���A������I���jʒ�pD�.��?_�Dϗ)��?�����J�葷+0!b����\�NW�d�%�e��@�x3��8�jiJ���wB����H��'xbg!���&�Iz�BAÞd�^aZ��!��B��
)���k���$�,s���*��w	JFa�j�c��H��!3 n>z�1Q��O��=�%��PQ��-&h��]��s��1oncۻv+��hq���QS'i$}%�><�&m���ᓓ֧�6��u&`���ů���զ�N�C8� 6���9>�D=(��<HP�c��9]�ss�&ep�(\v�{9���xԈn�eX��P�e��<Kq4C��ľM���z?8u\�)~p���u��i�Z�L���w�	b�5�.Cg�o �d6"3�e9�@�1�=>�\/�8O�h��}�5���ae3/�Z��P����Y���4�3�a�]b̭��u���^p�|��
o]��򩸚!*EY/ʨ�2,�\���W�I��zN݃�7�#�#�\ ���A�p+���+x� �6����o��&J�\��b��XT�Y���womW���ӱ(s6�����'�w)c�z��>��n�v��G�n�5��ƃ��d޿$#ґ�7�G����߫�b��AK&Ѣ��)�Ên�'�{G��:|��mvZN���̺���Śm�LH!sP+���q5=JeV	��-R��I�[�k3v�3��ɩ�}c�ʿ{�e��UY�3��&��~�]ZA�xj�G�T_�Ԉm��-��ԑ���T����G�j�	���N.�b\OX�19^�M�Ψ.\�1��D�Q��1��� �����_�6I��ɗg���;V6g�0n� u�3�˺����g��g���5���#>	�<q6Ƚͽ�*@7c�'g�-�)ޑ��	�P��3/
�i=���OE�vm�"��<YEF״v����7��E���u�&�V]�7�����.��'ؼ�Ndm��.oPH`Q��z�f�3�������J�L0�#�/"{����j��E)����q�R���#��\�������aG-�1(|? q艗�83���Y=��J��nc?����}Kke�u"�"�=s n�m����]��8o5ϯi�=!�M7,Y"Kɮ�[1�.-�DM@�4	ٷ7�?V�Yoڊ)Ák.:��JNP�ʛ�]e�wǹ�*���b��j_�=�:�6�wxT=�߾����8�w�'>͘��0j����3^�=���?~�ˉ�濄<��҈��fת�������/�(P
������j��mu�X7�<��~y�݌�~��+eud���?��Ulܧ5>����ab�s�[�����Ű�-=s*Gp���(�����W:x�Ȥ��:�ȷ�����)�|%E���`N�溄F�A����p�n��u}��3�y�����?ܸ������Y9���Q�6��z���I&5`�����~]}�'9u�Y�b!�b�l���p�B  �1LrO.�J�`(�O�]~�c�T��NH*�?��b�'s�/r�C*��8b43��
X|�����Ri���?����`�v+(��a��dD����Я�ɱ��"�h�����e?l�5+�7�~��:�&~[�}���c?=�! �U׋��4{�V���[�J��8����2��J�s�~#�K'�ǶK5�S��yD�: Սik���N�")���BS(\)�`DP���� ��^�!v�J�F��L�Yw/6s_��W���d�v�������S�Vs�ě�����z���[��M���Ȯ��ZX����dh+����a��J8�EҼȝ�0���}�Y�<����c �l�0����J��S]���}x>��ŋ�Qq�ý�|6	��m�?���a}�jo�HbE	KM���d���)�)����A��𰨄�DW���-|�2��e�^���8�"���������u�-�W 	�Jl�֗�@�ЭE��S폴��԰�Dj���&��g��#��<G��p�'���QJzzD����-���T��0P,���{veǅ�B��w���,���`*ɴ�d�gR��D��""^�˷g,���ۿƬ��Y�?�&���X����N�櫪�f����Pb�\�H�m�����=���Mį�a@e��nk�L�}�8Wt�陙m�\tO��� ��}�rż�22������;ʿB�dB�_�v+�4�N�Y��Ztc�����8�J�R^p�֐52^���(l\Í�m��4@��a���<o�MC)7��t�P3QU)H��P�)o� �"�.٩�#/}J��U
��(75����X��Qk�{��|̍�Ua�ճ�1,���a�������o]r�6u�(�(���J����&��g�p������C�ܫ�p�٨���K?�6X�Xg�K���ކ{K��P'�:A�]*`�e^2�o��"?��y&7{������/%h��!���z�uO��6'}��|<�ќφ�dێ?U��r-o�T�T���{�tIO�'#��ΰ��JG�V�ҟ��$ ��6+s|*�i/�ź+�C*���	��cզ����s<���?[�p���¯Q������+>��g�(�%g������D�1��G�Cz���� �V;i��@��ص.�¾v�\���2H�g�!Q뚻6ߛ�]-3/�:K�t�֒�&۲��9EmPd0#�V}}M�� �Z1�&���&�Nn~�m��
c�
����`�t���G�R�����J!��O�7ZL)���$���k"}Q��l�[>5�$��F�����~k�L��bv��N�{v�@����2I�� e٤)�po�/t��6��&�]ӽ���EZR*R[p

���ڪ|�p�X��� ckt����@��}b>���D����� �m�CF9�bz0S&r�嵲Ϟ��G=>�,�� H�,!���`��YkJ�"G#�tP?ReǼ�����N`m'|�:?^�;�N� 6����a��ֲtn�@���׹3�0ux����c�-�7��K�f{6�]��tZ�z�6�a�yh)�j���
�r�M��41���i�̝G*��3-|����G�~::o��5��5� Au��_�?�z�I����z$���X�ބ;����k�w�������5��28���EC��V5{����},P��YOר9�c*���� ?�;,���{�b���|r�����1h�����Cw&k�Y�|}��!�5���r�1��>�֏u�{�L�G*���=B������nӦ��q� K6��ѝ������L��($d��GwY3I\�ګ��i\D>��ٝ����c�NW+��$�8��!Q�K��)�H��(�_a�.��������@�D�@���MI?�yE�c�l<o��s?�������l	S�W2m��7y��O5ao���[��4�YO�A��R��fj��T�Lz��^����]��lI��2�*�5��ơ�3���O�b�.Kt6����!5�=���nC��S�=[K+���GK�^)�a�0���K&e]ŦB�8gqTF���'ڊـ���~��9]�N�^�n���A�G�D>�.�(Ŭ���k�b�Rbd��k?���#��-6� ,���v]�'5��]5˕
Sgʁ};�+�)����lm�� �t��5~��a-��WέI�cՒ7���#�����1 ۖN*s��dg柮*�2��JH�-�B=�a�0�,������Ж#cclL�9��;+Bj�ُ��[T�X;I��7�93_3���кT��$≘�������F1x'E�\��a(��fa������3b���]8����7T��^�&'=τ^�,������Mc(i$7���1���}}*d���?��z�tc�n�V^s4�6_y�;:��e�nζ�]�����{[A3�؅�W�������x.*��FO��bb��"y��1�zN
��cƧýC��<|eo��7v3�W�"�7��B���(c�����#VǅMr$��=å�d������P����=R&��Whڙ�Ɲ���54�W~I��x�8��N[a|hE��H���|X �a�:��� O�Q��&<�l���(���A��Xx�Xۥ�h4�ӛ$��ο4[���>�~�.l���D?�V�*@��ȓR��G�U�&:����4�SQ��|	�l龑H��$b����ܦŎU�1�:]���D���}[�s 푸�z��Ց��ΜO̔��b���l���V��4�jY��J4��	6<)�HO�6�fiF�;�]��{�qD!����b�k���$��V<��#�@/(��Ry��Tw#���a�Y�<�/�͵��`���Rm��6�ɹne�hOC�32�z�*���~��\v4qd�N_�+)��.ϗ�+�n#x ���R�~�nl�ya�9h����Y;j�u����/0�Ð6"��m�5�e�% ��ju�K��`u[��E����ӚR�?�S�x@�ж�j�7E�î�[̴&8o�l��ğ�]d�q]W���\*���|#o�xULQi�z�b|�	&8�g�;R@<�*&�1d���#!���4��Y�f� }�d��V'o�'�3����p�$
��H�Q9]��܂{�/D5��3vnZ�����S~�Uu7l����ݥ<��=p�y����&d�6TX�]�U�a�Z5�kDǏ*�2H�ˆrT�X��_~RU��݆64�ĭFa��1bx���?oF~ra)�w�f�
��^��7��N>��p��ek1�IOΎ�[��W̤e���uP����n2�Q-�0�hI��C�|�B���w�u��SU�[i��M�sA	,�n���
��\=�xp���m�ez\�Q����������p·��2�"O,TPM�9��k|"w��T4<����g׉'6�Pw<�`�s��X��B=@��oa��_�J�
���M��*ٜ^hV��X�_�<�&��=@�h(�4UJ1�"%�W������l��(�6F�T�z�u���ul�-Ro�Q�Z4&�4��:m�GR�QT,��`+��_D���(�U�Ԉ.��|���׾0��nk�&�	�MG�w-r�b��{�P
�𓘫!�E��39xR�q�n�^��~���	p�ُ-y����B��jM����D�í2��ޡZ�?��c��I�
�2����H�C�#N~'��q+��é��ɑz�%e�-)��%�����?
�mMQq���+P+��Ƚ+!� 7l��ڪ�М�F�o2RP���;})dE˳����)��)	�M%%���n+UĆτ�[���d2V&���ZB�B1�Iب�V��]�H���Z�^�V� ����'^b�q��pH:�1���4�rY�"6����0NO9k]�Gh.#O{Pr��b
C�x�ф�	R�"��U�'k[Y�_��y��'��gz��?�֪"�.Qȹ���|pM�`J2gڴ��,���A���k�'eM��ڃ��¿�'4Ĭ�3��p������1��/w�zڌۃ��[���B�H�U��N��2�)�ΈR���Ř���&��]%���&�E�+�cܨ�T��,��=l�h�\E����O���a���o��M͜���Qȕgc!�ii��\D���m+�D��W� ���{x��k6T�/�n��/	VνЦ�}ƍ�K���8�_2�q�E�� ��F]D
k�h���A��L`��t����N"$�6�tG��r%�K%��h�U�gP�4CE��H]C%{x�_�)��{E�'8f���l�	i�twl~����O����Mi�M�7�'1����U	2v�}�q�`'s���\����Wu�������@����uB�a������S���������*��<n�:��QʨLӱW@a�0�e}�Wε�	��j���#���z}��Y>��d��Q)���E+B'�������5���W�4�N�������j4}� ߦ�X��3�eѹT�����"�e4K|GɑM^z�L���Ja��jڟ�
7 7�g�.�È�G���ޡ?<w�67�ہt��D�l�Y�ߥ�$�U�,2�v~���_w�#��g��t���uA��ߟ�L6��Y�Yu�N[?Ω~!6��)�u<�r���n\��<*�2����u
$%�=y��4����3�i��=����;�f<N���SO�L�����͌B%���Ƣ��|�p����I]_���k�	���jw���;k˒�'������>9�Q���-�7�<�G�0�w_�w��*�u2j�Ƈx4�c3!�����H�T�`*�������L�C/$��>�c�Hn_;`��?�@s<�1a$r�L��UU���uF>W7����;;��p����t�\�,���-�u�'�zU�����k����y�/K6�Eμ~0�Uw�dnmܚ�4����IR!�������/���@RC����L��3-&w ����G�L�V������p�Mޯ��Oe2�dg�`�Ϻz�v q�[��|��U?�u���������Ǝ�oZqh)qY1�.��p}O����  �;3�ŏ$=��;9eC�=zw�YU��ԔbD����]�;^zt�p��%�˹A�mo�H���r�y��6���v���o�{��)nX�y���o��&G$�&�<��o���S� �@��0p��m��Q�K�	h�f���{8���2�I�������W#�E#�A[���$V�1��A���`�
;��`�BDU?ۦc��C�*jO=ʬ/��x��������T!�q���L��N�G��s"yB둻&�Z�e94.0k���Is0�쉏�:RGˑ++��@��Tp��(dR����� ��C�|���EA��_޹C����T?T�Q�a�}O�h|E:Z?���J)#��,��i��'2����2��;�ˣ�_������f�0_�.BfQL������[`k0Z��Ͻ��N=�J���;��B���'��W���ݽ��ҥP>j�rX��=t��Ü�[��H��J^�n/�c��K87�|�<,����S�C��7� J�r��|%��S -�HD��r�
l �$�/����qײ���ޘiP`��ԋ��xk���YjWԣd���c�ݗ��_'��\��O��������N�r��O�9�=�%�~���]�I��X�_�`��%�ߦ?�'�_Φu�y����n�󩚒�q0�`�%k�cņc̋y8��]���μ�/��P�!3�\�u�C�ydol,��B��Z�C8�du;�[;Ox�|�9����<���M�[�<N��8�Ɉ
��NZ�͞��WX(�EZl���e�� j��q��S����#7��[ackwR�)��ɉ�⤺�R̋�<p���:6;���]JS8l�`3����]�-.*Ä�2~L��~vW�l��
WQ�D+�jO��F�ޜP���j���b�E���6�!k�j�am�Q�GLX&A&��Nk6k����R<�I�},�R�֏m��Z�8`ڐ��)Lθ�??���p����n�Ӂ/<<| A?G@Z˅P�~
n"/�(�e����5`CEn�!��
\ֻ�w���Sm���
�Ԝi�J��������2	��W�%J�ox!a�%���"�����J����d~�D������yv��L��"�2G%�{Ώ(����I/�� Tjo�v��{05w�G���Ų�?0'�(M�Q�Yg����h�;B�z�U)<'�g�����fh}�l��	BI�Q��ٱZ�vG�����ez�7<I��eJh�(��̂��۪߫���u�sk���0Lʈ��0�"��H)<a�A� �j��妫.����>�X懶�ctN'�xFw�+}�F3b]�v���˵�������*Y�D�5ԏx�kJޞ�}���^���"����<��'K��Dm�_��|X�۶��&u0�F��销FP�����`S�����&��)2U�o�]���]�2���Z/�	,-���,}	�����ή�]�D^'~�bŹ�V^XAG��K��H�Gb�/�)&�q|܆| �'ߵ�QZ� Ќ�@��ɵKG�F=��ʈr�������e�n=!g�5|�-d?_F�(#�=�f$-;��S�U�-�mk5}d��;=33��~X���9^�g����` �>��~�\���>;m39��������~Ɉ�2B�'�S��n�م"{ӹ��l+���\��=-���sl��!/��3�}���i�?+�#�s�q�n����+[�}��4����~7t}�"� ��o�۳D�鈲m뜷��Pw�c軕�U_��h
�����7eg��#��֠#���A�(B\M�E�z�%??��d��xc<9lΐ�Y����V0Q��;#�.��a��Ą�T���9#F�d;k���-���qx- #��3c��Յ�ݕ��pgn�>����)A�V���N���h�na��*�Y�sz�(�l]2��k(p�
���� .?d��Ҿ�N-��8�ɨ	�F�i����c�1��)4{1�S��b���S�"�KNuy��x�%��Zg�;n�2Wj���{h���ou1�s�B�^~U��\�\v,U�.Bakf�0F+���X]�/|�y�� ��% ��@���'b+�ք�d���{�&���%�(ڭ���M��q���;���k
x����*+��:tY��Z'�3���KAp��:��y>��f����1媬�dQ�%��Ţ�L鈘2�a�
ݷf}RuV�)z���/���EX����]�x�VGMR���I��ӂ�ŋ�T�>l�(8ld�w�a�5`�?����Wy^'�VW�Dk7��d�6oX�Lb�9�U;Vi�e���1���#F��nו�6�뿅8F:^6|DՐ�O�)+�>>>N#��(����S�N�͓=%�����n�rP��O�,&s�}�|�zX�+Ǯ������'K�&vM�k�U�D�,��g�_f��^*ړ�f\ppE�L�^�u�e> ��v[2����&��� ���j�,<)w�k��d֥�����7�Ӧ���ʉ'�zv����v���4ut�U^V]y����uUbMw3��]�1�o��߳�۵�Owv���ςܷ�����j���'�k�b�� �:W,�̉P�6I�eֶ:X��\�mjz�q���oKPi�����C�K/#R�Q`�P�(�,�3����ta�`>�3�d�c��P�\JPwi'�d1>����[^��߫�"��3��F�~���#���_�cR艡N9P���4j�}�?#�W���12�/�A3��Mo�e�_����\�7l����jl��re������NXfd�"��>�zcJ����@S۬�.Y:r�c�1��d�OX��ti-;���@q��Ϧ>�鋬Ei��z/?Lfp"x�F��_���7��C!	�нp��)��!�֙L=e�O�wS%%%2!�IcWX�Uݨ�g�����?!Kg�<s# 43�1[!�A�mԖ�o�F�m4%
v!�3����G��C�+u�����!�U^;$�C9Zl�Q�[�r@hB<E�Uw偪n��
�*�Z��F��\\V��M�%s�2e5/%&�LT���A˸I��n��TI;� �,/3$���]=�skJ���a�Z����8�ߑ�4�-J��%�BT�%CQjCB�|��g{cx��Hl��c<	ӌHvT���F������O)&Y�/c�υ���af󀤿��=����W����ɋ*X4uy�Xj����D�Ogܷ��{��7���CM�N\��I	��e Ϝ�A�hO[p�P��ڿ�T	r��堋�	ܻ�<b�=�/$��- �H:�����ݍ��T��$���F�;ل�~�%돲i��E�?|�nh��o������7��uT�zq�$n�h��@���H�E[��]���ft���ag�����c�&��%��t{�n_��gܒ���2mْ�x:��#FG�(��=�����|	� ������${	y[���!�Jd�>��S�Ѝ��W�Ǘ�'�V����ޟ�P��8'(���#����4p����h�b�h𝖨����}�+j�ϙ����t�����K���u}�g����59qW�Y��Lj����d��_�Eo�Ǳ���ֵ��n�OK{7��A�j�+�^�ࡘ�Ԃ���QV�Ek@��:=�u���;2*	�]m���H�P=�i~Ɔ���* ,X�D����Ҵŝ{b�JJ�����(��G����r��6��̙�sq�T�3�R�e绩)�j����\��7���Kag�3�q����\��8�\n�dc�f�NH[�S&�!>����B帹����8b�����@�)�<�VYL���)N�{�H�T�SN ��ty����Q�ҩ���M
�ThEe!{I(���_�r�a�⇇�_�fwQ�bq.S"��w�K6�"E���~��]��b1%�-
hqM8��tĶ����W�Pl�4\��-_?Vi���)͵��5���;}Ж��2rv�kKk<����j�$f��E�dT�R#s�(���V=�^�t,ǧB�b�ۜY_OFZ��n�Ӽ+q���B��Ƕ3엙�2�w�С�[}D���O!�«zIBÎjvl��F8Z+х�����EosTO�G+�xGR��h�D�bАz�?�DgvI!�	��Ӈ��OhѤ���f���kg��"���`Ǜ!��h�Di���d�,�N �X��:5Z���_�X<E��y�Nۦ���������R.Q���UZ(%9��p�^��щ��Yþ�P2�[��=v�Pӿ�����k��ͅUg��j�KnW@�Uu�⒟nU����}�Y���<��]�J��9�a���9�V�ޕ���~,_Q�bRpN�_	9v��������}��2}י��Yj΍��H�>�&b!]`��'h��@�'l.PAe����[*�D��[�Ǉwps�\{*b��0X�Q}��7]m�F&�t'��m��i�2�ֲ��[�l��;i���HS��FD��/>�/I�cҫuޘIn.��,��M+�m*Q7Y�x������E(�L(3������̘<��`���Uړ7.!�~����ƙn���i�y-��52���+r�
�fB*U�djrܳ�PrR���;��ø�:�c���C@E�
d�������a���J,����=��T�f�ˍ;/���k1���
Ӣ���3,�����Z���ND6������aZ��CfEJ�?{I�s���m���#cx#����yJ��b���=�^f��͋�������`�ɳ�_��?��ޝǔ&�
��˝ۯ�"�t(<!xB?�no�a9�t�J},F�8w�3�"�ş&�w1�����;��q���xt���=$��|΢���})��2�<�55�������(��ЛWK(�>����%ѫ�y�'�9�L�I��'�a�~��SU������M��x���z��Q�g��.D"Z��#+�4���]@�&�,'�h�.i�Y�_9�$�͇�i��ͼEݣ�u�ε0H�����S�n���M�\�+Њ�b{�D?T�~_I���<����]*�mO�X��滎~yz,�t8ð���e$p`�k�	x���O\N� �[\69���}��S�b�t`ēi�޺��������fš��L��\[5-� I6���*��]$����o4V@
U�F��*H�Tz%B�N�uL��my�g0��}�n�k9�t~[��f�kb0H��x�5�:�n��
̇�j����3�

���Rh��l�oF��4�0��u"���w�Jn3�wE�a�B=��7�����`�%]�	�>����D��q��YC �¿��(kQZ�O���2�mwx�O3�ʉ��X.�t�"�����>���y�!l�������G�L~v��c�A�˨�B���ƖyI�Vsz���A�m�ū����]������$��
��I�=KiE�U�m/j_�3.v#��(싆�4��r>^6zQ���(�Gpఠ�>��\3����p��K��~3�i�[u�H�Q�.�	�o�I�����Uku ��
�T�`9�P��:�n�B.qO̡���`�`�Ui���ԃl���<�0�i}�c[��A�3k`ap�]����O�q��t�����?�f�걩+�Hq���%}\���X�����x��
 �I���!�8�E��NH�(���|2���{�|��Ҳ���b:C�l���vt�%"��!'�[*��c��ޱ��S��`�wg�y�'Z��O�5mS�-�LVݣ����j<���k��$2�yCxm9P~P�\�8�)�+e��{B9(x��c~+��汯s�_g��˄���1J��A���CQ�!�_������}�㒛��s�d��~;P{�(��[d��`FC��λ�������	^�Zq�|��q��*�5o��_2���&��6�wQ�kk����ڥ:H9å�+�9�ׯ�j��8����E��U7��c�_�BeaO��������<�@��r^?��|,��Ը=<"<=|������O��O���՝�����-�Q),�¾��1�*��F�9�+�#�r򒑤<��S��l��X�󺍁©����n�S��F��K��⼱�v;�!�F��{��>�=�;��6���=���V�NL������Ȃ��%sF�����'%h%��.���Q��	�zt�T�����}�H�%���JIi]��t��_L��bPn����{8����Nhm�0�P�%'����j�H,�$:�`�E�L'jͣ��QYb�5:��1�J�ɨ!r�/���v�E�6�E*�����;��pS�Gh��,l�L�$�9�:�~��F���l`3��@�Y��2�6�.�f�$������-\A��ȥu9�Hs�򀬲`����J3�����D���7�&�a"�,�j��
� ����맪4��Vf���J�$��}�	�OzfU�F!SI��j���ף6��􂱴.Sof�NS���j�����}���9Vv�4X`�Qh�8v_t��hy�J�B�����p�mohak�>�fz#��n�����<��:�7� e��i�Վq]��X�9�z$X�36%����r�G������˩��q�$�Sf��)�.��F�ө��4|x��6�^R���E�a�6[��X��8���Sx�w��h�s ��:��H����[5��Q��4�^��!�k;��v���J�C�������~����#P��\��#<���vc�\j�.[Zu���l��2�ׇP��S?U?�o���ܷ��ޟKnƖ�m�r=�ȔM�~���ֳ�+��>�ܭ�� ڵ)�C$C��fc�:����g-����/d�If��NB%�zHfrC�7f-��hW��Bb2//��kGC��9)�Pd��/�\�dS�*���v�*r�}��Mq��zX����ě!pv}V��ཟ. Vs���ѽ�B�h�(��씎�a%o/�L�R @M�q`}��k�ZU��=9;P�/o�+����fR��\�4�D�g��|@#�|� E\�OpIf��Jj����d'Ľ�7p	4�����XW��ƽ�J	I���^pH�7��:b�b6���s{G�UoFGG B�v�s�!�sn����������L�4�K��5�Ob����5qa�s���2����'(��*挖4�q���u��ڻ�_x꼖F��D1}��a˱��)�KA�����8��i_�S� 敚E:�,�γ��n½`�fAw�����찧���#x��3����"T�ڴ�L�+�|Qo�)͞��7&��Q�%��~6�GlرFO<��<:
`�:T�����x�=+߹�vQ���z��V�T g��;�\�:[��@���Jz�n�}O�&���dV��>o�����Bk8�_�Il�ۘ#�/n ����wVd�͑�֯�����M�)�
�9�=c�k��4`���A'����jڄl��W[7�\������f�	�PwΈ�@���T>-O��x�奚�C/��3Z4����e)Z"��ByR�h��<���&��?je����Ye�n�*φ�j=)"�`��>�I��0i�M��%R��b܉�,MC��e2Vw]�K��;�kNN�ղ���?�B���yH�[�L�f����&�=:��!!(0�T�����^>u~�|��0IG��_����(D�8�ֿ��n�͙6��c��!x�2�"���Z/�a!�yh
���}
�΂c�:J����J$J(ϱ�V�v�d9��I��[��,d�?��1��/��-\�ϭ_�'�X�M���|E��_MyDʂ�� )�i�̙����#(��R���ֿ���+�����2����V�m�#RF�fU�l�ń7�@n5!փF5�UAe���#�&�#��&ۦ��Q{��0���&(�ݿ�(�)X*����W���NR����y�e�Qڔ�Mp�o*�]���pio�ۓ��~wK�."�z�9����EZ��a����F� @�D�R-����O�O}���N��]	8��H�Q��h�9<O�զ��0[=�yU��tx�*i�B�!�b�%!��W�&�"�72���T!o�0��3��]0�X&�b���G���  Blr�tEE5��
�p�D��	�*L��U䛰�%Q��=�]y�?�t�Z��zz�(�C$���t�.x��'�ίɈڦ���ֹ����G��'u����7KF��D<��)��'5��a��8HU�S�!��(�dx���n.%��q��)፞�ɤ��
Wܷŷ��1)��i˵6�9�_w��������*�BA��/���DC/b��`�#nY��M��ꏚw/�n�b�e����r���Y�����,?�J,	�߼Y���:T ��3#�z�
���EM���3�piDx���5<�(dx�;�"T0��H�3�A�q�}
�#Z����������pQ,��*ܽ�e�I�o����ʨ��`�����;'�3Xpw���m��w����%8��m�7��k���u8�S]��z���i�[>�+CQ '������� c�w�FF�$P"1�?W���$.����`b*��ю�a1���v�?0$g�J���a���1m�إ�0��Q�IP/
h�s���{aBd�K�W5̓7�n+U�%6�W�F�CgM�#v���'�w^��@��"8�P�h�g#hxAu��^JFw���Gj�Z�:�!F
��I^��[(�����	���Iˍ�Z��0�nzi��t\���vrJ]�!x��cP�^��/����з3S>J�8�(�Y�����2k���#'�n0g(�J��[a��։窗�^c���u�����'=_b; �LB���\��c
k�Y�kg�~�q�5��(�ŧY�����8�
_��Vsl�پ��뮥��ǫ=�/�FY�ղ�˲��}�@�|����^ۼ�f%! ��^y���Cņ(����I��b��FC����XBm�l�@k�?�A4��c}_5q�� ge�+ ��-f�&��:l&�|g�87
��'��Y?�m�Կ��>t$j�����-���,���`�5��k�e� -�>>P�>J���ڳ�S��We�,��+eg�������_��<����T��D��OhpzD����U�X�Z�z�j��f� ��/����r�X4n}��H�8k��MV�yzV�ð�TI=���x[����&�̕�����]�.2�b:��<��Az��>�]�ͯW8���=^�Gj�ϫ�tq�$B������6փ��H�	@��N>�u�G�`)�>��p[P�&�Zʆ�/e�~\���q2�����j5J��ˑ�/Sz�.\@MӢ�k�)+�Ҥ�e���.�a�*��|����t��o�2��q'����KWr*��݉T^�u�
��@}թEI��#���<������T��]��v?U�+�֜�Q�D:+�w,�21���U�V%2��X5j--�Y���ҍ#�Dve��������������	����f{2f�S�.[�{X7Z�h7���7:�$���`��Ch/���Qߍ��t��s�=�.0Y�[ P����Ks:���G<�Y��s������ b�o5�0����Ep��݅������ J�D[��<�O=�=�|�5Y1�'�_�����0Tg�M6 [�Y0�]����tW>}x��Y��������l�і��Vˋ��I�>s>vV/�D�wG�/Uݧ�A˓֒��˓2m	�y�\��K��5�4��H	.����;����D+���sf���4UEV�y�#�O d�:�l�n#8�d�<�W�!��4�P�D��m96i����
��|�@��?�����I�����|�ח����dK^����5��P���kn������4�֓��#B���s,�z��P!0�N���3��q���L�=v*\Y���}�w���=JnwqÆ}�h��,��.d��zE�\|Ӆir3��|���de� -��'9���	XSӽ^�&���ŹmU.�@A?�����ϟ���^]��vË��6�mv
C�O�OA"���[~K+.�T~��̍�����\ �YX�R�p��8�}��@P�]
�b����
ٟ�__~ɼ\*t'��1�m�Ęȟzlo��_a�
6���G�-�6�$��}0�ܩZ�.I:�{���؄��c��F���N�M�G*f'E�`�Pi&�dM�<bLV����h�?8������!,��]g�N�%wI�1A_t�1�����*W�\�My���P>��W^�m��71[��@��Vӝp9�z�Çhژ�}瘃�QvC��^���4��]]<�c��s�5����������m��z8�{#����|�Y`�e������ /���ib���t}�cBN��+��t�S�ÊJ���_8��R�F<0Ҳ���B0�XJ$Z��>���w~�\�F��>54|��9�U�pZ�;{�5,��H"SQm�w@)�UT��������߫��7"�+�7;�c|哘4-�f�� �3 ����^i�j�I�^���Jx��S�x�v���A��V���:�*�ز���C1�芵����U��\f!kmF�_)���W�e��d�S���n�ݭI����|~���0{$�^�
��`���ʹt�7���}3��c���U���OM�oP���������������mt�z�����]�Z���~up\�.J��4*YϘT_�Bv@)��x~к�̃�S�E�w���Ц̓^EL�!���UC���bn^r�w��ʚ�{���2����=;��n7��O����܆m���Ɍ�O�*�©�ێv.�m�q6���3S�E~)�Y3�%m��n��U�߼���D��|[����٣�׏(eg	�t���Nbe�<�J�d�ߵ;�x!_]�]XfHZ�`���&�dBLh P8S˪N;|�6��tG�Q�-��y���jǮ߫V�����$I6���h����(��~Y%e���T7r�@��|V�0(�ų���V���]����	��J���/c���)��Z�Dv��(d�w�{�Rǃ������F<NN��Fn�u��
S�ڇf�w�%gs3;��(�U]E[�Xa�� >��Ou��cLFȣl�:�DC���(J��W��ɅQm�̀k�dQݻ���Av�W\eJ%�_�)1Bf�:�����j6s��i�G����Pr�&u	f"˷1Ҧ��`�Rks�U�Q��h~x�m�4�0bjg�]�Ql��l>p�#�d�%/�G~�{��ʢ��崢z�H+6ߙ�����.|���<Q-?�:���2���x j	��1}�h����5+I�8�$n�~w6�{.|Z��s�Y˿V�+�%|m�E��2��[���dq���D����fL��,�l�R˅��S��#�׃W@��m>��h"Y�$��P�� �E$���ov��X���N��42u�u5'y+q	�g�K	�B���b/��͡��A,4��BT�iA���x��!ֻ���$f^ޟ?�7�$2*[�.�Lz����q#���Q�t+v?�C�b1�z�����(�q;�A/���	�n�2�晴A������k8��H���y�l��.�΍ů3��t�*Px뉖A�D�.{^=����G�A%Q��#1��ϸunp�KbQ���N�㽍����̉?���T�3F��i0���	fO7V�Tv�s�w=�f&������c7�틯�`Xz�d���%Z��yAP����WJ��+N�` h���{�t��n�3�X�]����Z�Sҡ.[��B~���i�K��TӍ8�x��yO��hL�j��}-�����A�e�������wz��5�UL>_�ΙGx��zq�yM�4�ɿ��91�?(�NZ���_|�k�K�$V`|T�S����a�x�C�t����q&qi-@\�fݺ$#�����<��}w�(�y&|�
6�5=5�w�7�]^+�|f���{g�n����Z�4�8�l�e������#�ōbP�3�CI�"O|Ż��A�VG[��;ߒ��C��`�j����!��k�>Y�s-��.�.sc��/��R�#dlZ���3�w���ߴ3ւ}�]<�
ġ�]ᔍ)������CE����8�<Z�/C��,��B���^���-�ҋ�j�qy�pOd���k��:3\��"J�t����t�X�u+�r��P��<�Q���S_��%�pV�e#�G^Ek�8(�_���%.�7����t\�{O�'=z�����j��L�}��Z�n�9DV5e7$��CJES0r2�T|'n͚Zs�^�����Ħ�	=�	W��e�����.:�{���L����Ra���=i�Ǩ}�A^-�HC�S�@�5�AG�g�[˺ν�D���m_����=+�i�۟�\�an�/�b`��1�L��%>Jݕ�*�Tj<�j��_�SP�G2yu���7_�*x�c�H���>���Ӭ���	�Vu+��D ���n)$��4D1o�sw)�7��ҹ�$&��/�|��E�hyX�IG	�FFe۹M=*���s�@�d�뾘���%H�n�?�T�p�^=mn���I�.��<d\��<,��&��>.ΒB���_�Q{�<4�l�X�t���;�|?�7���#+#G̫5�N���(�&��%��g���ٷA$H�>�
!缁�1zZgFْ�. �	�R'�B�k��8̹�#����V�4i�����(�O�2����5��C�U^�8��
��G�����h�yJ]-�#��bJ��F���nL�
��N��Vv�MF��p&�M�(J�h`�1-�q*���#`�����<�6缭/
�T���F��Gb� ��&��9^�3z�g��G��&m'>���L�V�Ӝ�i���K����K�A?	����9y[.[��u�f$
�W�3�|9�<$NaIK��$��T�<rד�'��,���3^�'n�y���J�Z��ld1_�E�j�5���܁�=��K?��4! �xH���<a�Z�wBs^�=���QB�Z��1I���f�zo�U�Vw7*����gjԐ��ʆ�s��T�\?=�C!��8��Ї�
���8�������[N$�(��F$B�UQ��c�w��'�e>÷K�����œRM; ��O���-���Oz۹͵Zթ�:���#��en*�EZ�����ļ�.���� ��	����K 'e��ƶ�̘���צ��ء�S��$�D#�e�{��<�R �@�7�ޑ2V�t�]M������/=",���.�_{����4��w�����驕sn����j��ڽ2iPy�ė�=�Ϸk���$Pu�CT.�!H<�����^hB$I��r�Yt�xl8[��3s��od����X58��|���<g�R�;��X�
�)m�� `;�ܽ��-��lT_��E�1��q^�܇̳y�2C�`�08���x�[�% x��矉н�D`�\E !��lJ�k��� E�5�Kګ��6r�H_���o�:J.#���e˞�p�<>N��Q�Gb�ɐz�:�>�)ĺ�I���b���◮�u7x�H2n�Un-$���Wi�	p{�0���_W��y��b>��.�8_��}WD�f�����<��.0���U3
,{��X�=�?�E�u7M��J)�ZÎ�Tׂw����]p�C�Hd���S�g�kcu�@�u�
�ǘܨ�DXy_�#�"����#"b�q��A��vq^���շ$c<zo��VqT5���wm?�+�����N�.�>b_�����B�$��h=t;漺pu�(&����o���s�u׹}��HG���Y��G�P�/�s�I*�,��Z>%��p�@���;��qk,1M�N4W��:8~�iB�0��@�����/�/���������5GOh�|
�k���:� 6�͑�{b*k�ν�,໶��s~��^�3D����2�`R/*�A/Z�?9F*��*��*}l�ҭ�5�����}���W�G4�vE&RÝev�IJF��?��@��ǁ�Js)�g��� ��­�������2�155�_^����NMb�S|MՀ�{O��M���W{��k8�ɠ����n����l��;�n,��3޾�1�
��;T�����wt�(�n�ʎt��O���H��h'|0#9wD����f�� ڏ�/Vv<�����Y��ާ��W�*�2��'��^&�)���Jx�=���N��4���x��IZ���]��>��;,+�7�2jeD�`(��07���G�MTt-�M��#���ׇ�;�H�f�c�4z`���tI�����v��#n�I_��/��K`��~�s��d'�\��AP����b���j*y�鷀���n�4�R����$��\��
]��^�2ݬ���{Օ�؟�0JfN<�����C��f�	)�k�ɢ��x�� �����[��,Q�)�p�h����')j�;�l��31=07K�5O\�\���-�	��%YI)�M���l����z'���l�s� t�MMX�v�̐�<a���L)����]i@8-x�ZA:"��JX N�d�����!o���`l��b���X��_K�Ą2@�g��/���A��+�XYB~>*���8���;�b�?KҵLZ�q���?�	��ꮶ�W,�J�%�d���4KO_N���)��.fՋI$����n� JՕ��0T�d�;��W����n�Q��e�7��ŚHw��H��O�7؇)���ꏰ�jw�ۘ��ӡ�>L�nsQ"�FA�Ê�����$��9l҂��NaB�0�= $2�с�<���p){'���J��(fnm�������d�5}�e�|�~��Bd�xb��6��ѥ���R�
��̘�^�W�a��W��/����]��.DB0X��� ������H�I��N�Ő�@^�]p�Lfx�=J3�C��+�NS"`ߩ���R���T�rȳ��0/�/��DJH�_�U=��$ G�̹����?X���D$�l_�r�@e��`��j�Ji<�	i�UluHI��|��%�t
�Lݖ�J� ~;"���e��"KLN��'��CTu�u|	�o���pd'l}���8�|��� �7�ܿX8���
C \���fu^"����+ �X�!�ݩw��ey����B ^��Wp-g�6��[�ȟ__db(�r����m��::h���:�n�<�vxĜ-����e|���L�E{+X�۞Ɍ��3���J*��b�Ƭ^��I��5�~�&�K�ss��I?7;ҊP������+�լ��p�0\0�3kz����?��g�Zx���F����g9�+�͇V�DP��q"�k�g�d�t���@�P_h���P�e�#�(kL����2zذ���Ը�����|<��3�1�tf�$�78��󼨷���J*��0����e!����l�K+�JɱɃÓ���'��[��/V��������!��[x@�xX$��O����Q��ݼ{��Б�K-�^�u��dd¨��Դ[�h�+���j�o#���0�D4D���SvG��ؽ!�1?Fw���
kڥk�p��I[�'a����O�W�1�Ę^�s
�΢6�\s��hr�3��΃N��
��͓v�VA��-�@���Q˳�&.wGt��P��U@�;Ǩ�1����ŝoq�H;SՖة��n�j����w��Jm�@��~D�O���>���_H0����}�Vv�5�0����L�	6bF*�L]8M�+#�T��u4��8_��A�!b/�u]����@�6�@�����-�1��d3��]E�T���b�d�C�_���;�>*���t����\z٣���,d���j�f��@c���B�|������RK��@�oP�`R���`�ʰb�����<+H��e�P[���*��f��%{18�M�V7B�Чx\֤y�Q��ZZ.�;�ԌRB�F��w�U�$�0��AZ���.���,|9�B�|��� �ҜI����J�ё,k�?�	䶁������վXN���nհyI��������4/����JA��.�&��z��~]�$����� �E�_�H^pϙ�e��^��䷾p��Q��1��\ �p���$:�m2xa�0t�&�K�1�X� S��'Vo�"�L7!��t�Ie��q��V�}��u�Z��ѵ���o�`M�S�U��@��r�(�����@�)	 ���|����ߠCm]�<�>x�U��)�\I�3	��Yi�wTྏ�<�Xìqq�t�+�����yL����Z�����F�R32T��+��>��!�R8�o�y���Y#�G"J�Y���^�B?4S��mmQ�݁4��}ZtC���S0CH��f�F�[Ưx�+�"��i��wcO$��\��.���iwj�2�M\����yi�Y˩D_�9w.ʱŎ�
Г��yL�e�(d�6���@���2���-���e,��?�������#��F�3.�Y���S�<UI� ������/�;�������n�<�~( �w�u�GW�{�i�����%�c^%a�m_eг�<)f�q�R N�J���*�_��0��fp^�S����U��� U���Z�D���JH���EQ�����j�Y����c5�����5�D�*_3��y׷a��#��?���״bn�bH%7���B�ʄ�u�}<H�4ij5}ͻ��@m��`h�e�@��q ۸�]ٿ��0lB�E�Az9"/�;�7�ݚ���� �<.�s�%�^������KZ߄U�PRv�_�ۼKU���Gʇܲ�3�j�Թu'c�'���-Ӑ�,�ߩ��L�l�	��m)�[�\�`��y���,�I.�T6�/���uU�@;tC?�en?C�[��9P�@n�+��ő��,��������SP5����W�uv��&���d��Z�B�缌̱�c�Z)l��1ãz�J6k���t��	�����/"�	���͹�j+�8y�s]#�k��.oz��g��!��g/�eп��4F�rmxz�V�K!�{{ghMǇ̙���ӎ�Q��b��2I����4�䅘6�@Ե'z�sT�Z=�[@���>��I��	��c~��8#܂����/v��b$�s�6LG�"���z;<'f9�Y"ե��P�\���ӻ'��8�m�:P�>�������о��ι�Zv��i���V� E�dKr���x4��X�4,���,_\F�L젠��X��n�Q*$������x��`�.�?��tV�-�n:@G�1v�|�����|D��7o�$/o����$E�+w�=��n�v
������.'30.�50;ND�}�O�7����'Fj�>nb��Jh3��� ��"�D��)�	ҿ���Y�啧������:#!/Q��~��g���0�5Y�39H~��W,Hf�*ȝ����9P�͊!�MM9'� ܃�8�?_�o���6.9�XrN�Z55�Ʒ	7U,Vz%�d:��x�M�mRw�w�k++��f;^!ưhuVR�8��|�d�FY�`#|����!��������9��f�~q����nͻy�T�o�B!W�u2�e���꒐	p �翐�J���_1o%�9h��"	b��zs+��;OJy�^D�%8s?t��Q<�}�J�h�bp��Z��(��[�b��������Ɗ=�xºG���˃��)Nz���U�_��ߵ��Z�۲)��/��DL����Α��>wkW�55s�./L�~Α\ϣ�X�ƞ�;t��!���CB$��J�|�|�٥L$�(Hj�/���~�.�K�B��Zp����|RT�� {j�"��Z��H"���d,�Vu?b�ϔS�\zUB�U?�ɦ'���s_�x6��zw�H�v-ށ$n�ކ���J؃�fKO���Jt�r��n���U�i�����r��JҖ��>"��47�^�U��q�~��d�{�Ó�K���:�����ȋY�7̐�ſ�G�h��G<��8�3��ʻ=��롪fGFN���W��h���z�p)2�Ϟ��_~�w[<Y/7���#~!úU��k:�I�8��n^1Դ/8~�a�z� �;�{(�8����.�$����#w�4;��w�����"8�E�䗮k�Z�0_�l��s���_0�TA��@>oQt.�ΐER�r�5�Բ�®ܴ�Oۻ�3��-ܴ�4�W�?&�8��qW������,�o<�O�	zG��5��������m��~^��3������^�>l�F1/
�|���\c�$TC�i�ß�2�t��ߎ��b_xE~��5x�t�R�ة��W\�l0.a{�ԝ�w����Y<��#��cʿ��+$.	]b��.G�^>j1(�K	�����	��rm?T���ZjCaau���� Q}�c�� 1�����l�Y,� �����r��M������K�T.�g,T"��тIzv����<����;��ϸsng���o��w�#2��0�Ǒ c���,����܉׵��sLQ��^�aK��뻟��
��U�k+9������*�q'U�[�&�>���jml�W���Iv��E
J]{��S��Vj� d�0_��J�ѥ�\����_fs����mWE@��Å9K��/7��I�%�sԫT$��Ex���rHgFI�b4�s<�$�����?'��>������ݘGϷL&��o*PS]�����G<]l�DS4�����(�J�6?]V�Z�Dl*w��OW��ξ�x�vŕ#���(w>�_�p?|��{\<�	���@"���q5�5!�|�v~�EY�XE�|�.GG�!��^��i/�mP�Q��8m��^��n=O�)���x.5,����D���z/2l�r$�����}៊��:������gE�~TcM�_�oFm�=~�	�D
�G�^�7	�/J6��;��� 0��
��S�<�r4*h)�gc�H�B��|���lU%�����=rT  ֨"����.��d 4���[�H��1�4�TM�J(�իzArp
�wp��yNo���M6�]Y�&��b�k.E�)�hFs�%_�D�6���uE����Q���\�����+Z����)t%T�mX����tb:Y9�;b�>$Aч����U֮8����Mu�m4j�@Z�K>��.�O͙������' �%��?�˽�/zo�s�? �F�T�.ʃQC�T	�֫�ڭ�g��fA����K�2W��u���)�4�M]K�[bD�ۓ����!�L�/�]�u������ӈG�RT��������w�n��(�HM�/���*��a���&��7L����0�A	��a)Dگ�:����ЕD7e��n����6.�0�6�
���{�Ol�7���d��@��L-�:H�<<��+�
nʷ����1w��2�N73��\��ZJ��6���;��+��r���b�=�	i��g�8��������-��g�
p��UW#e7����vR��- ��%�N��|��L5�/l��3��t4��U�](�?�<�{�h\�{�|����f��9��T|Mb<yj�O�㾤�b�0._��kِxc�J�K���|H�����2���*�&s��IO�"��?k"���1��٭��䈵�yV���M&|�!��SB�j���_��IoHp�dg�ڿ�����
��jy=��n�T?GE��G�D��Y0N?,z���Q֓��{�&0^{9����,*�_30�A�h�^�h��R�J|p{ot�����{B��?BlrXm'f�]'���]�Ŧ�b0�$�G���U�[��׃��x���:�fB�W_�6u��[7$d��\7<��`'y\�#�_���-9{SG㈒
�:���ln���U�������>����
�@Xȍ�G�_��
�?�IE>B��f2fe�K�un_P:H�V�HW�ى��Gv�+X�H�:a]Ye��5�̥D�ivq���%�����CCAi^�:�����oA����G�g;6/���z�%��e�Z������ç�7y%���l����[�G1�b�`�����Ýx23á��+��PzKߖ��J�W�\z�=�W���4��	���Rk�I��;�++�Z'������Vj�	#O}�&�H�,�V����my|��G�2�|�����j�n"s�v:e��u|�θ�7��1%�O=���QP�}���t	��(Y�.*� OW[�����Գ���=�x�IeN� �N�p\懍��A|�%?�������d�@�b6s���4����ʖ#oi����y�6��J��� X�g�z���<��wf,VV���!)��x0��g;�1�-������Ij�c�l�_��!��]����P���*!��5Z&�԰R+�0k��?�)�޺̈́��b��b(���UÔ�8GS��Y!��ٓʥ�]�C�9"5��ͼ���٧��ʪ�ӡ���Y�ɓ�,�2x1�80��|��j��'�[����}z��t�U�7��:#]�{�s���q��������I;i��� ��h�4���HHF���'^��z�A�I�������ώ �7'f�$�'8<�c�
�s��ɟ�ѭ���ߗä����Jev��r���>hz��j��G6i��$�>;�<�n8��%��u�K�hd�[pb����� r0mG�����Cb�����'��4�]A7� |� ����&2 @��	�־�a=�6���LˌQ�"|�vD
�nM[�NI�}���ٖ��v���N���}�7%=##�LnaS�3��������'288t��9xPZ��׼�%��ޓ����C�ӓ7�i��e7I����Ai��Y�󞲰�A��י���8�>=3��-���Z�<~����}�c�q,�b���r���p^8� ��ye����*O�Si��2������13�ADs��ԁ�����1T ӵ�@,w�_Ȧ(��e�	:��㨢e��EOO���f�6g]��7����2��$�-�x��6���xl!�tzq.,,(��,�`����W���C����&x�*6�²t� �7�U�i�#fҮ�1~��"|��l���dAS�֖nk�#�;�������c #�_�cΚ��d�����F�M�ϲf���V��Yw\�5��K�b'�mlt`������ē[����w3��Wx���H�BG�QA#�1�
�ST �.2�b41w���>��g�:JG�"���/��>ϗ��oQ8�4�%āf�K����&�'0ڭNfC�A)_07��:X�g�D�L�.p406a��&��A�E2%v�1����F��-� ��u�D{�-ANn���:��Ɵ�ȌG�9eka[���^%"M�p��JP2�`"���TkQj�,�� ԼOf��Rս�d�h�5� �ͩQ�i()�Sdjl�S��,����e#S�+|9I������_q Nr��Qf��E4�&�}�_?l� �L=�Ji�_ɵ�K}��=<��$���m^����k���?/���`��9��%�?���� Z�1 bM`�+e/)�z���Ҷ��$��^����H� ��P� ����u*�ThLg  8C��|���Iއ��u����Oo���(&��"�)�������}�Q,ȣ���LFЋ��$��^=�.�*+l1[���,��H`� ����7�^�_�P�Ђ��N)S&�g��:+� z�_���t�<�V�����I ��ȁG.\\t����3�����_$\�Q�J!�o ˰�u��Rz�Q o��!ṴX�թ�x@C[X���1$�i��Rd2���D����,���Y ������e.��'ب_��/@�g��O�wr��}�ѹ<����\Ǎ +5=/�ұ�	}�ʫ�_f��eFZ���?B;�����/P�i�ct���w��֫�>V~���?l��3x��Qh���/xhVta���1���b�z���D��y��\A�U���z)qo��ۿs�u�0�-�#T��Ҽɉ�
ɱA�T��G�Þ�1��a ;aˁ�O��y�y����_�j�{�ǠΉ�rsSё���X��|�t�,u�x'�"�=�8��.�O3�]��;^a8㬦���p"�(GI����}�+ա�trQ$�1��;*5 �Ob)}�����A��?�QzN��v�3�:׈m�S�����(�w\�Rb�ڨ0�*�#2�Sn�u ��c(h�������[��Y�l3�Sx�7K>�<;��I�\}��c�3D# �J��0�^� �,cF�8Go��B����.W�ğp�������kҍ���^��K����|/FL����6��q�ߘ&��%�������2>Z~��:�.z��ɿ0�� �;%~*�ka�bW|���Gf�3�0J�\�������#u�p�N���ic��a����L� �"V^rKn�u�dU�Շ^�����փ��泲��.��� 䐰g*Q����;5�F����uB��%C�3��A5:��N��~s؊%]��X4�'8j�{s�	�IsGͥ��V�93DAq6b1  ?bx�c�W�5<�w�<>��;�d{���P=a�3Gd�R���W���`��e5�)��+*^{��n+��(�N���D�f�H$)a���,��!A�Bg�?Qx���_��,o�j���)C}<���=��b*ڔ2'���4X�L�û��{>�a%
퐰�����D!j�9ؑ/�ذaB,�Dh�b�_^����:H�-<�L���v"�t��?��Q��<�~�_N���M���� -"�ȁ� /x��}=t�H^��t�c�Z6u���X�\�R�?�~�ry�	N'c�pC�Q�=}@�89B�v&�/@���k�}C�?c�cױ�AR�vN�m��2���Ԇ	�?s�,�ԓ���+w5@�̩�}�A��T�ߦGŋw�jw��;��d�S��É������1���$��F�0�ɹ�P��b��U%�a�/z���+���  .n���dо��]��l�����m � �9 �g_j��)�)�q^��J=��CL�$`eE�	�q��S`�Pa��!�L��{�:r\5����.��xO2}����z!z���*7l��1�=�����s�%����6�ԇ�� �>(og�c�U� ��>b������\�b
�=.��}?5�J����7}Zڧ�����|:�2���ԾO�,'d�H����و���50FB��l\�b�.a[��u�r�eO���=��P�X^O�M�3؞�"�$�;>����@�wʧr���#�?�t�S���>\��8�����$��tj���Io�3���8�j�JK��G�m��(� ��a�����*�)����m���'��<e�M���{�K�X�i=���:$4G�9�ƴ�X9	k��^,�-�MS�xs�����+q��	P�d�nb%��{2��{�x<�V��5�ۗӵ+�/ hS�E*�ZZ7F�H�;�(x�|����1��!1�9��}�R��ǮKGں֬�A�d�@2���,e
��7��NQB�D�O���*	d��u�a��_ʅ�E��� b� 8�*xFЮ>�3��'�l`���pH!���$R"� ����六�'�8:�OԆ��#޿~}%ɇc�wW�FI�|ɭ(��-~Uo�s���.+@��� �+ɒ�'�1gi������މ�wib��ҏ�L��?�iǓP�������7��6�7n_ƒbV��H��	�N�<�y��+�I���7�b�7�s@�z��׳�Z�!L�� s�<s$ �D����)�<	*+���8�o���@]��V�;2����f�� ;��o�0NU^��'7B�ⴔ�z�mQ��ӗF�h}��1G���>!��^ �j�9e�S��z ��o��d�O�E�[h��K 3U������d�×"x�]���:��i"�ғ�f��WN5�j� [+P�ʊ�Qt��d��� �#7?�I<������rsa�db�`��c�@S�⨄ku��&g��΁��'�-�]JׅWb�W8�$��ơ>���Z�s	���A2��/�����������	��,��dSK�^�5Ϝ�9���30���8$�F��\%�G&���&g�$4�H"]w�������Ɠu�{��E+[I��� ��yB)�c����-�ols`����ö��<1bì�+�])��]x_�+��� ��F����Ť�V�7Ev��:O�&��%��!	��$�)]��E'��)���uK���ɋ�[�ς b�~��U���1�x��8�aD ʒ����w!�%8μ��EqT:��#�P7D�l�T�}����i�8�L�eF{�� =��kn��o�ZI�e2Y�"�:0)�/m+� 3����h�1 ��-Sa���NJ�Φ3݈T�6�R�X� 2�R&}f<��1
��q���}];�8�"��Gq]GM�d���49,��e^���P�*%��TBN�_�(�X�v��ʰ<&4���G��4? <�~����<�JW�x9̒��s�����@�9A�$�k�9H�����f`t �ЗH0n�9+ T�\p*�M�"L;�גG$@�3,Q����Xa]0	��Oa�+z��NlXg��;5zj)���c�~ޱ�=�գ��A��l34��Z�E��=XG�8���w��N�E�Ϭ����m�]/������3�a_BI�+S�(�����<��q���YV��RRI�'�M� F���PI���P@VR��#2螵���Ҭc$�0��F"����Y^Yp9XMC h䚽����c�W/�[�G�݅�`(1�bs�wJ�0��c����(֯�ȬF�-+zP��m��;��e��Τ�a�+���cUF�x���4_4����BC+8��H���~ Z��=HB"m[��
[���(���ڒ������4��e�S-E%z鑩�L�0/�?�\w\߲߄ �&���" ��4	���E��@D�tB�+�P��" MPz�*U��k@頂���}�����|����=;gf��wf�9��{E6��/��6��/�]���s[�����t}_�B�T	T��m�Ȯ<_��/:+Iu�m>��u�W�!2f6��I�7�m������8�.�g�W�>����Ș&ϫo/��)�u��qq�%�L�g�����	C���S��8Fe��b��NG�dƩ@e�8?"���(�>������[�&��)\[�����?��,(K, �$L�v��k�˔�����ŀ��}a���(礑��b3OC����«�vl���{YB��P$Wz��׊��a��
U6��|Ӧ�,Y�D^�~�%U�}���(��|��$����6itY�N�/|��[��=�|?�0>@f��Ѷ�=�;f�w&˛��D
܍��韋kx�%�a0o��� "V�9j�[>m MU�i���W>���2�(��]����܃DJMO��0/����@@X�r3��-t��X&��ia�U�l��<�^@K��,�q�ۭ����Y�0G�/[W�������G���>�k�71� ��B�#<��E��3"r��v��2�Z���z 57�)�I�}e{��[EK|W^�F�(��y�c���B�T�*��~��v(�Tf�Uo|�fz����SǽMI-�^�p��T���|��)��0 X���	o-ڈr8�U��Ƚ���I�����O��TM�%��`!�ԉ�t�n`�6j^�T��J.O�sn�O���{�"˩�L����|�̤�H��/�:��\4�خ������&��OT���&P���˒�6�ٺ(�3�4;�@�t�	7�q?Z�6k�4}���V���M���$��t�*�L��`CS �Q���M�΁)�O{h^a�oa;�g)���q�e/�aL�� o#W��u��S\�0i��5��� ����!�U��u"w���ůwLt�ty��i�T������ɕ��UR,4��'irRU�������#��:��ܒȐ�����W��g<'�������[����Ӥ���F�'� �4�p����~�!���n��|Ţ��N�~[9G�_|0��Ǵ�wh�2!zy4C�AA�`Q�:��(����
Q~�r���l
�o��eu�����/C/���+���*�=I��}��#���o���ݓ#�E�5���
L2����lM��� ��=<Z�	��k���-�ƧbL�p��o8�����g���ߡ�=�p+��9ղ/��%���(����?�O�]�Fl� ��e����l|[�����*W}���!h���Lĸ�(��W�,�%Y�����u�tp41C���B=f I��f����%���۷o+��f�*u��'�����&A�N�Y�Q�)!�����G�u���j�O�J��}��x���
�:����F,]֓�T0���@ Xj-C���t��s̟�*3ͦU�io��Hn��K�q��q��e�x��t�H�y�*R��/3�0h�x �G�[�<���*�@ï=���B�����+Qt#!_���8��ee5��j=��ֹ!�~��L�"�H�1�ԋ�����^���c��ʧa95�E���|�ApL�bKe���	a֤�+���eg�}�K�Rwʋ��d,qXz��c�C�[r���Ka:k,0�_dm�\��
n�[�����,;��CJ��[�k3�]��Hң����~��5��	K�/�^J�=ܪt���^{�ٳݯ�-n��5=d�ĵ�-}y�j0t�ZԮ�*X�]KWӾ�W1����х�uU4���cc}���Q��9�NR]iN|�(С�T�/����Rk�Y��q\�2��=`垠=�2f���D9M�9 ���$XY�p��ہ��RFC9�Fm�۶e�n�ҰZ�K|`D�ѹ8�~&��H�oPR,y��Ch���Ҡ}�;����-_��wo�zp���ng>�i�侒ͱ[u�ulj�߬��a#gӮ��ت@Z.tr� VA!UP���57o�g��g.�*F���c���о9��y��/-ʲ�q��A܅Ӣ�:�Ę�X��Y)S�I�R��������g_W����h)�	v��h��D�;��ɚb�]�w�ӹ�=*k�ߋ��aP2����Dy����$~���a����T���.��Ԗ�'d�~t�����W��>��3f'}OS����<�� !U]3]���zhKT�J��04�v�o��3����-�?ʽ��$��2�,aؿ|�X�2�Z��^l_p��[D��&
4=[�������d�[���?�7J(&qt3��+����o��XMу!����?�tHxoY��ȃi�W0�r��'ұH����м
�M�z�=���2L>	[�4��}s,+|\�I[]�[�*��h�:��`0X��G��".U9[��b����̦-����
��oJ�4}r�Q*�ݙ`U�����ќ
�oj7�|���9���ZY����@��qƭ͎;@�$�j@r���+�?~�6�
2[x��X
�s�}۠sk�=�"�	���*&>�U��kzuѾ�6p���Yl��x����,����>�g�E�
�M�N�Z�{�������}x<�xrMԬ*���LY�ҫ��������0^y���N�J�ޣU�bR�>�
�b�����t�t��72���DV��g K��Ed 6����uA���;���R��t��_�Q�3?�N��ԥ��M9�C���k�Ʌ��@������¼��Հ���tWP�P)����/LhkkS@4��-A��w6wd}�w$.#� ��
-�L=������0+[0׵��{��͹�<�dl,~����������s0�|��n�rX�'1҅?<��nsm��)�R^��z����=\��j�F8O�t��d�;1�=(����F;�h2���@GK��5������Y�{���ѫ���G�*�_�$;C��Ս�N"�YO��
0l�@�ض?�P��3k�{����	v4U��f੼9�`	X�"����Rߺw?	�ڝE_�*�>�X^��7������'���B�X��*�<$)��O�-������]H�Z]�[Z|�
���ft��� �� �<��qd!�����*��6CQ�o2+��a�5vt��p� ex�o/��}.�)�LT�X;w��5�����]�y�o����K�r�A %d��@�/��L!L#�u�Vs���eE��L$���I���w�c�W�*���f��c��@�9s�\8�M�9�k_EPɇ���:ۥ�_.��hI�Ϋƶ,ә[."t<��R�'e���q�jɴ%��aؾ�H&<yᕢ���s��[��iWdB^�L�~##���]c��8��i��Φ�;���K��ev���Y݄�o3Yd�J����@z��ͳ~l@�p){��,,-ͫ��YT\L	4��4�_cǤ$��ks9���&�IW.��W�ĠwdY@���Jɳ��7�����j�`xR&z��O<?kB�}��\ȶ#&qwt����y�M�QH<h�ؾE�}+�e|�*�iPzb��:�2�g�C������_� �8�;���U�����2���k���.�+}vt3���S��)��{�ZY|yp��wI=���S`��J���XTQ�xm���X:j�������0����_^�)4�|�`g)���9�-�tgz�]�,���Tm�Q���e���5�_�[�{mLjh:�G��,�E�Z���b�]!���4Bq�����K��H4al��p
4�G��8���H�������u�U�)��D˰�Z�!���Xdݺݸ�"�$=��#��u�W�F/����F�r�D[��M��0�;��4�Yd��Y+��*AZX��n����3�S��������$�����r�prO���& G=��k.��l�V��|�5�Ԯ��w�ߟC��1����0��]��7���'W���g�uk�*������
4f��Z���/�����`H;�u)�B��47�$D����ܱh�G=С 1�z�W�;r�����Ȇ=Z=1��^���C�lK���S�f3Ǘ�_ɢ����05�i�H�U��F�|_����$��}ƌ(���k�0��|��z��q�+ߍ�V��­�Pq�����~|g�ڡ ��G�8į�l�f_����Q��Iɓ�)�S��׀~"Z�<�ڏS���ɓ+U��4ws���njo���,��c�&�{�W��1xH!�Ʊ&�����TB����MO��Ό�z��\��e�t<,�P #��x�l;��7jcq'���y����3�ym[C(�~y�)����!�x�S$�?�l�\dlB���Y�o���NEw�?�j�п�1��U�$�G������e�y� ��.y�u��Z��'�mk(���s������Ʊ�(.��75�T����i���%c�Ю����*�d�TޟX�̜�G6�����L�7;����A������8j�Wr"W�O���$�1�<OU�:eTQ��|^�f?�����6�[�
<$�;FFC�D���e�uO���+���־ko;�>E���H��m��!eh���c�c������5���� \��sc�����H��B*{Xy0�MA�N:��k�����*������6����1�Z�S�f}8��j���i塸:0p���*�}���'���E`�+�?�6 x'-�*`%�TP� pr�FHpA�C�X�tiX/h�go�W��Qy�@d�����OM$3���v�d$h� ��}�3:�M��=D
��9 ������/�?���R(���#���ЂMԲ�Q@V��	B�d(���<��O�L�ξ�P~����3x�Y8x�� T��c?��r�=,(|������Y,5'x>��@�졈�o��x��	��ʌ��: H~zh#�
W�"������%�=S��
ݙ|��,���\9{܊��Jfx���6$��E���݀���yk8�?Ӑ�p��C���L�z�p�gC	J��S��ɯ��9]d^�1� Y�{�<k�>�����!h������\��!zl*�WO�ϓ�SXl��	�ߊϡZjz�o����PK   �a7YN�v4	� m� /   images/4949577a-1080-4c93-a0f7-9bc81c12f32a.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   :Y�'���U  �U  /   images/79f1f6d5-8698-44f6-90ff-b688d5ed2669.png V@���PNG

   IHDR   d   �   b܉{   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  UMIDATx��}x���ْ�{#$����+v����z��P�]�a��{A��bGADA�@�=!���ޓ����̞�d��BPr�����Yvfμsz{ߵ�װ�6���T>���d>���G ���e4�Q��j>~���5_����67��	ai������� ����������vt�� �W2�S����|L#7a  r��0ANmG���4�	��C��Z���L6&D��J�� a����FA&�A�csP��������NN�� �Z\��i"�1�����L�����X�b�	2$�x#۟	0(����Sjx��7	A��a���]A�E�<�\���'������?���K'�5,z����_�_�)���7�Q��J�h$?7A���)�*�V����jj��YF��A|L�)���U�^6��n���G�fdQjX5Y�N���>����Q��2:.-��0Afm�MKb�#��K3�7?+�D�Sr�?�DPB�E��Qp��l69�ںF'��4Sae3�5��D����jr3���c�uTc�-�3zo��Q�"���[��S��
:*5�r��軬Z�+Iλqs��R�(L�Q��L�`ѻx����-*z�f��r�0��wٽ諭}ξ�C~dBL ��NG�顔�D��ڴ0��]�G@\�4.jlvQym�7R��ZZ����m�����x�>G���<��:�W���	j�k8M�C_7|a"~�a 5�:3e=�՗�)} �q=�<��������k��F�g?.��b���rV���j����n��e!�"�蘡Qt���th�0�����p�)uP}��8�!V�?��J��@EU-�dK5}����.���f�0�=�R��Of��Y#4��6��q���Y�G9�3�!`|��C�	G��I��_^5�L��_��U��J1�@H��h�:�����O�-�]>69��;�UD�Տc�9�	s
"B��7�w,)Л�}Qp+ssbB ]rT]06�z'���w���ڗ�q������d��FE҄�Q�]�H��QB��Z@��{�~�S�ل&Fe\�g�O-k���H���G~��%b$������z����^3T6�>nAz����a3��T�N��k��,��~�/7�EQa]0���k���|͍/���7=���*n��ul̶WDvh�E�0�"#�����c�>ة��Au�F�=���`��h;�}v
]qL�;��^��Oe�Mb��� �t~w��B�B\w�K����Ɯ���ugu(%��W&�2v�ίh��q�*|1�8f榥y)ʰ��4p8���y1���7s�B)�椬�zy��������3���O����m��G@�Y����^\yP;Ĉz�qΑ	��T� ����=!,�)��&�ElH��t���p�_�?<Rs�Y)t��q�����"& �Uc��x��2+�fZ�_�=ӟ�I�EI}M��Q�-7��0p^M(E4�	ǚ��/p���.� ���,�����g5�yT@Û�5ad���۟m�R��X�N�QQ;�æ�$�c�8��4��X
��c�O�OB\ =zq/:��h��#��n�*��������(**��;w
⛛��������)44����(==����(<<��'6�MMr������=�l��5}�Q1tׇY��՘��*ґ��>ޥ�Mf��,Sz���o{�ܗ1��i�Q9�=Bkެl�?�5ʹ�1p�g&q� �P�8����`�Y4��5�d8�I�iw�_~�&���L�g����@	��XETc܈(z��ޔ�Sm'�	����/����i���x�bZ�`UUUQEE566R`` 544�u�����'D0` ��ۗ;�0?~<���l�ev�x���h�3�d�n(���6����U�M�!�$xG�+4���>�[��~�3����f�9΁�\�BcA�0-D���U���P��7����#ɗ��.����Q�̱[���rc:��8鲓��ы�ȟ߫#b Y@,�<w�\�1c-\��JJJ<*J�b �AAAr��1�ÀĬ]��V�XA�~��H�رc��Σq��Qpp�Л0�Ja[��-��Or���
(-��s^f��qVZ�n`[�����L�u,UC�k����`�ǁ PWH� ��h�aI�Z}���}>=��)���,�l��Iڵ�C�H��h�Ѡ;�Mc]݃�[���jw?$H�ꫯ��ߦ�+WRmm-EDD���H�-//�;�k���D�������BBB�p�����?з�~KC��o��N:�$y.$�<��yl�q=�OV{�<��Ŭ��qYv�.�+�*��)����~��y�n�P�R�b��_	A��.�!���<�!���6��F�_\���\?"ӱ�0�֘<s.5�=�Ѥ	)���B^)\�C-=��C���)H���jH΃���f�0����R#�����^|�y��ęam޼����
!���N#G��� �gs�~zڰ�PZ���,�u��t.������	�G�~ggxV�=iq9�W�7�cۑ�ק�3���K��,H�	cGӰ=�����y�z��gEB`x���dH �4���������9 � ��!��p-��	��1�|Hޏ?�H���q�B H�{އ�k�:�����e��E����/.����b$��pʱH�ǂss� SY[��%7�N�ή�
h���CS�����S��ݺFJ�MeNJs�4SF��i��0�%�������.��o���P@��xp=��.>��wv�7,�E���{��iѢE��O����<D�H��E��U�u㒴���T�(Y��;��'�����B�uH���6���7h�\	"�_�Yہ�eS�b����x��C�Rr�=Qbh�P�ᴞ�t��%����Nf�w�3� ƦM���o�e˖	�a����h���'�\[�Ϫ�`3��TeFii�Ge),\.���������ϧW_}Ul�zoJ{`CG�DՕ��;vl9���LRH]7�!ze���lrH��&���|��8G@nqg3Z��|r%)H�p���kg�������6?/�f>3��� �.���ǆ��o	
��9��6?b�#�ƍ���/]=u��g �[\\,Hr*++%���
2aԨ�>� �-,(++����Jz��iԨQm�bH��F��@�U�߲9;�������7�� ����ި�soz�ƥ�bF�Н���<��)�n2�C�Ȇ�������h񹛍|�ؗO��	��,�����i�Ի�!�g���wPbH!q�N�����䩯[\��!#����x��m��%��^z��<�	b�����(p/l����pi�X�W�ciP��πc�Z���,H˶m����׿�6����4||jMM��7�n=�g�5:���2.��5�s���E	�;%v�	������pJ�K�8'SZ�C�
&���imI �Q��PV4�|Cl`=�ԭ�o�6i�9�U&���|fR���1�1�tp�7� /d�.7s�9b>���6����3����yH������믗�R���{�eD�vn:�i�f69îir:�6�qc���粆�@��	�[n2�m��k�^�&���T��/<��fI���&&Ʊ�O�cvQ]p�c�Nm~����=a3B��of�I����aG����í]�d�x8xy�����32��U3j3�Z@\p<�{p��竗��8������=��,H���/�u�V���E}�'0��C%��g�57�pڞ��˪ƀ���x�G����OtX\'�wuK�e|T���Op�tm�u�AB��'�o#� �����j�8s_{nb]Bp]8뿞��@��`.��;�"�����z�pc�x����P-xIE
����:D�kAD��ǂ0J ܋� jJ�5�PkfX &`� PI� T�|x�������'P]�I��{$mY�0�n�@L�����J�fܤ2n�<�eɀ���=]pLd�۷���36$VStF���Q���Q���j���L�m�]�N��6m��w�,�4�J ap�p� &�d1@8��yp8`�>|�q�UX@�@Jp�{��\@�G}Tra�{�n�8�̀��Pn�*&��)�qӯn��
8=�m�/Q\� 
 D���A��ȟ�+���S��1�[�S��j;%g̜#1G[xz��%;�ċ+A��P'-����b�gF��@����q:���;��k̰px��y\IB���/�Q].�C�=�Ў-��d�����D)m�VDj�C������|c.�ɯe���E���+�
u=x�l����e1���")� C;g��8����S�U�|oNwh:����J�8���{ ��5X@4����p*��;GaA=Bj`�/��BQ_���b&I:��������)>���oP�e�TE��5���{���iC�NamKA�
�끈a��Fcz�#Ж ��O>�D��*�.�i�`���kq�Z H 4� �{�2q^��
 c�a�&��+c@Ͱ0�L0�~x)i���Au���J��7z�_���(;�8D�������D8��H
�P]c�'�E������E���������������j3��8�q>�a�>�oX@��;oXZs�yi������:t�癠Kp ��c"iņ2���G/WӇ�3A:������`��v��Y�f	7��Rxq�0�p�&�=��:�os���&�<\.V' �`؁t�ă�x�8{����0TM�4p�A�1�x���)0�mV��KMy]&9\Էg0�Idc�l%^
����/�E�q�4�j��8j�[cU@��Ps ���8Dai���t<��1�!fX`���k�����t�m�y���g�� Z��F�W�ut� <�Q�`��&S��@�
E!�<8���!�z���*!�AB�k
]��r��u�R�VX ���́`g�p_G��a@���#��H�D���F��U[���@��Ȍ�v�A��� d��TāXu51���s�D�980��
oX�絑Aai�
�U��/����B����Bou���Kg�+�_R�T��/�t�RA$��Ѥ�Q=#ﲫ��$���p�zY�*_`�:<�j�e.+,�� U3�a��5kִ�!���}���o���jG�&!<ш?J��#���u����v��Psb.���2���q��,-��3,M�h�y0�C�fh��5� ,<�W�Z��0���'E�-
�QiU3�+E�H��P;E��$޴8��\�io����d�; �Ƶ��q�Z L3,mbPX@�ڟ=�BU� KEoX��&u�A�^�zy"M�mF��Qi�^Uv�/A"���&���?�F�ܚ�ut����f���Bu��q|o�����<��`��|^����Cn˃
F@ �!�ԨU	a�d��hq�uy�m�D���,�ЂH�9qʙ��5�pa@����նoX���$
כK�j34��W�½�K*Q�?��Z<�\��
+�+����>�.{Y���Ƶ�@�MZ��|��!��5�.��Z�̰`\����z 5c�i ��8Ĝ��PX $���+�z�[���2A����jt��|�������|��p���jP	�*, Mai
�#Xj3�a�������7,M�(,H�f�;V�_�+>��.����ƻ��]F�k���͟;*�btT����[��RpG%es���̍�d��)->m�ä�嚛Ҭ+8S#dp ���v�쮄�6C;E�s����M6�R��,���l0��:"�,rvm�k	bq{%�VaӀ���Q��]v5�p���+��6�\���C̭�澬=�R�5�,�T5�x6��]8�q�7���NyX,v���ߘ<�d�4�in
ÜqՈXcp�f\���j�ޚa��WX�z��zh8��R�5��gs�K��j�[���A,����no�Y[�5�p�sg��{vt-���Y��g����Ka������Ҡq������"�"��Nׁ$3HL��t�X�۟(�#p��C�������nj�DS�eWp��3,s��̩��`�K�8�A
�fx��ԉ9��s����.�d�e�5�W8O���C<߁ x�>}�Ȣ�����n��Oum��0�4�g���[IͰ4���pԧ�1���,z̘1�EE���xH�G��~���5�p��?%�(0���=�K�u����ns�>knJ�|g��nW����y��W=X沫��a�� ��XZ�Z�"�ށ���K���L�3?�Ġ�]�i�QC�c≉��0S��z����ԶRm�Q$j[�X�#Z�0�ҥnfX@��`���P �&T����r�"ARP�5����&VY=�äb��٬}�F|H���B�����A�  99Y:ȡ�4��]�UwS�����S�|G�ܫ������toX ���kv�;*�J�X�سg�v�#3��-<���6Y��/��B�2��R鞐S�3�<S��A����Z���E��p�UH����Ͱ���l����a�.e��qfX�r��V -�{����fP{h����,��還�ʲ[�nkMucRxU[㣎:J�����
��n7��;M��ZQ��:��DEFg�4Ů���,�Z������AG}t��	�ڄ9�٬�8�G��%	�����Ĵ��CS!�]v�,�Բ+�T�yH�6�A�h������b���u�Z��`��, �kw%܎`ib�#X`��/�X$G�V:�a��vi���2�DY��V� �-Q)�wg�u��7G�d.᪞��4�����fX��̰vW����c�,wk�FjzgI����SW��}'?���!K��趵tk6��6p�\{�m~jԕ��Z �C�@��4��TB��*Iai+)`i:~w�p=$\��B����`�"�q���K�kpP}Rr:\��X�,%��v���3g�i��*0��.vw�î�[u�8\��������O̰�<��g),�
ש��w��駟.s7��V�t` ��Njlv�(ᢏ�=�:'Ű1kq#XS`(a�L�"�A�>д��eW]���ZT����r0��*]�R3,�i����}Z��f ���&K���8�.��U��UNr6s�l��	�y����e͔��'��i���z������TY'���;i�C���q��J���nn%5/i3Â�0��.�ai9���Ao� 1@H�V�*��ܒ&�'��qE�/#��`���hlZ UT��գB��/u�1��c�=F�&M��T���W���U4ī4�^�&��0��̰��+~A ����H��s�p�	m솪*�1�q��+������*��D.g)���z9H�h+(���z@��?���ǜ~�,*>�[q̩v�sJ]�e�e>��|����W]uU;� ��^�C��=���YT��u���Jj�^�Ni�*#!!��=��� ����/�=�]��4uĀ3�eWݍA3����6���j�3X��0��'�ۺ	��֔q�:��YBv�H�u_G��]PK9eN
�W{�L܆���֡D��|�Ѓ�_�j��:Zvմwg%\�݀�%\s
]ai
���ӧN�*K׼�x�e��<����M�,=��l�1�D1��m}%�?"���+�MVS�VI:4�`)�ɓ'�FcZ*�}��Gm���Z��:쀶�`@B�\��6��<x�8�rH�X� �̩���¢"��]2�]_��R���B�dl_j,,��`{�� r��x)H�م�K"M��g����������,_ޗ��6����T�u�]'N�wZD��dtFQ����?�f�Xo4�uat� <����hG��,V[�(r�{�2�cQ̆
n�.&L����O�s���n@j3Tei���,H�w	L�IL��AH��竚��]����&�I[r��d?O���sԷ�����qqTR���$���`h$�k�.AT�v~��H�{�'�}�y��7o�����V�*\5�dM��y��- �B�	�#�86���������ɒ�z�c3
d5�Ŷ��
c������3~ͥ?�j�s� �wj7:�*@�Ð�U��Q�,�od��ٲ�oݺu��LW3Y���^�v�@Zt3؈c�=�N<�D٥T�|ޕ?]���;�ax[D%Ma���u�����0�A�=wAa-�ZVF��N��b
鴵S�����F��������\s�������0[�l��{a��e��a!9�V��K�H=z�h�,�{>�
��׾�N�Y��u��3��������5���?"����7�����NF\X�{}��"aW�� -e�S.Z�R��8��S=�F��3��s4��m4T%��B;�̼'b`���E��hz��?DK쏱��m���k�_�쑽� /��⽛��]� �k� 5c��5��b��Mn�-:�{4h՜�v�h����e�4�?������?ҁ��$��d���t�!c�ΑG�����\��n n��h����)���v4��@M��䠯�P8uuh
�%����9$�B隣_	[R_�DS��@�\;�/ZHCz�e1a�M(at��zT���6q�r�ΆJ��� ���!���7����b��Z>��05������ؿBX&m�_��̃�����i�ֵ4 #�{Y�TÏ��w�F��fOH=,��ɜh�W"�@ANA1:���&�Vo,#K�����N�1�|���}�p`S(g�.J��n-��Cm�y�t�kj'|1ξ؍��BJJI��;��ܗ[��/10��@u9�t�������d�UD)I	]^��y�Ų[��?�kWA!�Cb��L�>��{��Y����ϱ�eL�wL�.X����҅Ex�d��*�&k8�N�n�������0��� �'�6���ϯ�7oCs_FM�y���L�����@�@�eNn>5�EӠA��ǗQN^���_5�R�`�?_�YLWL_Ao�|0-X���7�Р>)d��wy��_1�R��D���)8:����O�=��6dU������	��,Z]B�?��޽mm�����Ө~��	��P�TSUI붗P����/4�&<��v��ˉ��DY�UI'߷�^�8�F<��/ZJ*�'{`ZZT*v�R^���8�(Z��H���.w��B��� 0��Mt�#��s�ѥ�K󗬣��iX�H���f���I��X�l���ژ[I1ɽ��c�ӳ_eћ�eI}�b�kxG�o%r^����7�O+�ˆPȀt�-a;�h@O�ߋ�����RiAR����UPK@>��.q�/��۫$%�7y֞�C^�#�U�+�Va�ӓ�?uUTU��U( +�z'QBl$��`�+��1������J�i{qQP�u$�lA��g[�y�=���� :��~�N�/�g¤��GL.���ٴ*3�bwɲ��$�Dr,�<���ם%f��$"��A�*o��ՎK�A��N��6z������Ԃ_��TЁ� �W�F���>k���9�x��T:l� *)��m9��fS1�e��`��Q`�]��٬�jѭ-�z�����7SU��j����B(&6���H��PZ����|���.��!����
�8��!`�=p��c��L����Ó�A}��梪�z*������/��%�NI":Erl6��*��J"�(4$��]�aG5��c>����JK�C6�J=u4�At�ĸk�e����ɜ�l�4&P�a�7%�z��Rb�?��e��o����3�ŕ��a[m��壚r��C�Q7#�yt;������[� �[v�Ж�j�l?���{�w���z���J��\b��e ZN=O��'���Kǿ��e����C�l߲���⃟���Q.��[b�����{��0ͫ�D���7�mG��^X':_T�^��0J���������(�%-kW-mɯ�#��v��I05[c?^��!���+�^��L@�����*�����l<w@Zm�UG��FR\D��m_�SE;���nEy?~˧�B�!~�ǆ2���T�0&��xk������D��7C��iCV�q/���[�\̅���]�������#S貧W\
3�����;�������;"�wq�c�h3�\�g�L�]���`?
b��/�^�a;=�lK]�n�ͯ���_x������tۛk�Y~��K�����33hқ�h-�G�"����;��{h�������S��Άx��:��#��O9TZ�L5;�IǍ���`�c���YY�.���K��!�=�V7?�ǥ'��C�GѶ�:z�]픘`���4ٕb��2Z���.`��7ҋ_gk�PW��FIQ�{�?./���@�A��]/ ��$�:��g�XK�2�O�@���0S���h��}n�&��G&�M|�2�A��F3r��KC?kp]~i{S6�/�^�~;I7��A���C���%��i��X���Lz���t0߿h�����.���r0��O�q�s�kkh�ٽ��'�S#~��rV%�|�0����U�� 56�w1Q�{g=����&��;��C���_�pj:�bf���|�e5�.5{�ۇ�����y>����X}�w��"����F�d㚗��.�_�"���J�u`�}ӄ�򹕔�����z�vP!�4�>�a��*flS^��=;)��U�6S%@�Ȍ�iE�3�X���=9�^�6��<>�c�
�GWY�,��#���"�EV_���;"��R���*v�k9��M\L �t�0a �s���`�f�3kk�i��*�z��??��&*�h)���^t��k�Ax��,+��nE�K�ElCJ*���C����N�Eg?���-�و�,Rf�6�^쭿x� 9�v����!K�X�����~��o���V�?rp���M�����V�\��<�rCn5��Mճ�	�d�4S��Ĩ@��k�o�[��Q�ݲBJ�g�f�JC�m8@x]B�x
�[�3���6ֿ7��A7�j,�{���4wU1�cd�wA?*c��d����x���%UM�3i9~��ƹ/�l�ߘ4R��>�D��@�MU�ts�HҢ�et	s��^O��f�G�|��c�-��ީ��g3��χ=�d;p��hz�QL�Z��g���Ig���ɼ�UXK�s��:H���,p�A0P{X�6�_ӖS��z�G�*���3�9��q����?�]R���r$q�0ְ�X�])�>��9������J��˥/��6�s������"o�[�� \7����5�BD���=ƪ((�[d����b� �-M���Vy\h���1K�#�"���i W�~6��3�Z��׿��Z��x�1|�����ݿ���9�������SȲ�6�����1A��B�k0KԦ��[D"�fw��J�u��<�<��1�S��,���^�W.y��v����]nf�r�5.�j65�ɾ�&f�`�݆ x��`��A6q9��g�: ��Qg��26��%����_/.�Y��ѧ�aP��Ki�#�S/|n��Hn�KY��3��ا{�XcY�v@���F��S�K6ۉ�G���y@b~a;X�N�ݬc����}���4�����z�h?�%��;7�-+�s[/��	53�m�O����2��d"u粎g�����jn{'���uPaQ����z���!6��9VA�m�) �ux�*�v�`���UƳ���� �ꄞ�Μt+;'�q�ԏ�x_?���zK���-�0��3{��s�3>���kKi`j(��F�q��p�"����,�]��Y*�~��N:���^�p���$j�+���w�������������(C��d����4ZǱ���wҶ|�1��� �vŶJ��r�Q���<����K����=��:aL�Ho5t4g��kߞ�E~<��N-�t��:� �1"!���{'�2'��@k-sr)��_��/���
䀐C8�8aD��"��t���Íb��=�� �7#��WV��7��lI������[^H�2��l����Pz�=���݆���&9:�&r�>�����mi*�g��I��yÛ:�%.t#K
l��}�0"wdvg�8A�ae��t���*)�	rb�����<!M�JH�o�J9�h��FgcϮ��:���EL���U�U�ji`s0s��e���Bܪ
��dV;���=�M6]pd2M��U�&�a�T��ğ��0v����|ԥ�i���#YαǯkJ�?۫ f�?�^��J��k7�3M�Y��w�@�Ds�G@��n-ڗ�52�[�2�c�xp{!)W��F�85��,B���f�� ��5L��X�}�z6*O`�d|�g� ��	w��x	�� �h�����'�I|�A1܅sx���8JG�x"�HL�@&����&�{b�؃Iv�Kw� 9_�nGZ����H6wG��;Xz
�L�ea�ST�y�֩�n� pK�l�ǆs1G�s�`�}�٫K����_����
7�ϫ��s��!�*�g�cG���~�����i3�e���q��HrEM3��6�Fg��Ż] �-���k���l/a�Z;���9L��WK�!�$��/|��P5.��\��/��j������?2�A�	�F�œLpi[rG�ps�zk���T�l&�l��=����/���MgO�-݆ m�\�a�B(�5�t�'nq73�9�����ax�h������y�9���u$݊ �O������۵#��ZSɛ�7G��47w�\aj�^��:�@�9�l6�7��nE��vOc_�r�a����Y�R�|��9�������B�_ 0�c�E��+�=��a}"�}]�N�7�=ĈdC}h�(���<�q��|�{��s���F�vT�?�N��,�7�g#��Q�A@���K���>�"����RV�Ɂ_�]v��cG�R0����#���/�J����=h �����3#���>GD/A�ck�e��m�^�΍Y�:CLЇ�`�J?�r�(��������2Ɂg������zg�����Ϸ������}��i�4}�m�t=��|��1WÓ���j��Qt=y�������o���(��%����RE� 5���M�\��/��Gj�������MŕM��oy�r[�h�ǌ��Y"Q��^X/�q�A���̭���:��P���#�NT1���@�*������8ŏt�[�݂ �I s{D�mf�&F����7�8�'�1�w43��vӣ��ТM�B��T\̞�(VOW��S���Í�3i����ޣ��sn7y��Z��9�#�O&�������b7���PA48}
��A���[@p�F���Ә0��:,��+p�r �έI~)d�u�.����\�T�P�������ۄ�.��N�q��ؖbz�]Yu�|]c�M�[]�BU�  ��J���=�i	-XcF��a1���H�]�-�8�'??��h}����p��,���AG���D�|���r,�[�R���:H� -���U���*%�*���v�Ev��Z`d#;��e�Q��"�&��9���ZI�!�pi�a�Z\@3�,��j
d�B>��a�4��|zB������d�E
\����w8`��a$�ɶ���\�".���b��3h�CqH�p�̮���t6�������Z:yTd�@�O,_,56�Frt�T��(7w	!A3�[���'
ܵ����[�bHk���9���^�fH�H;H���!h�Y�:-:h�Y���O1�&�����-��]#6p���N��T����K��Z���v��ң�mv�5��E�$�������=�qx���7��-��:� �#�_ĭ�t��{_�:{d��"\�I�����?a�C�S���{���<�ݬ]Y�"p MO���n���,K��Z���ܩi�w�+�[#���U:�A0�v��W��b�׮m"v|6=[%���ˎ�nG���G�!�D�NS���cU%�����R�j�.]
 �\�V��m9��%��b����.u���}�1|�mT�Ɠ�dZA�Z����(�I�t펻�T>[܄C���	��(�5L��9�@K(�b�?��cp�pv�#��s1G�T�g�y�9��Z��G	o�&v�3-s8��d8�~�ڡ���.�yc���v���% �kr����J�ꁋ�K��4Hd���rvՒ?�k4$���`�ǅ��3_l!����W_��n |(�!�Dk����Ȝ��ְ=�-�bvk^Y�(��v�g71:OTRQ*FQ,>2@�o1#%D"��֟�Ӈ玎����f���W��0�*z�	���L���1�M�%^� ��q��{��di�Gn
��e�+��aDF������#���Gz�7�ѿ��+�~)�B��?������������^t�|t{22�Qm�"K����k<�͟r��;G�4a�ě�s�W�z�Y���ޘ8\b"��*�W�l����O6KG�f��>�́���h���&�Gݥs1!2��8��M�;��X� �Qu�pYă5��5�X-��7����� �����okKDRjX�!�@:#��5�_�sA���]��ޜ_#�\ 	�}#��>˪s9����wfD�󧼵�����Ig�6�i�|���j���Gy���5Z�����\$9����ӻ��Y�%J���y�OF�z���+�\T0s4�����Q��Kˌ.v�A.�"]$�(GT�qԈ����vث�Cc%�|��kh3� CJ �����;�9��)F�Ҕ�r2��2<O��zD,-�DP��tb�P������T�u�Q^�?�/P��5 :���
��Yl�z�,�A�g�JZ��\^:�'gdl� ְ�p����H�3:�!������N�ggm����꩑?�D��w�b�ӡ��&}�������jN:Է�hT��t魂�ʨ�/D�3�#F��G�mF�>���I��a�A<v�w��DV� �?'d�.V��8rG��ff��<�f�x���#2�e�������R�:,Y�6
<%U��̗ۤN�ŎN��>G�9�3���>�(j݈@ـ @t:�!�,�eZXgWI�Fw}��SĪ���qՃF9
� �,5}�1/~�%����]"�H��b�&���R���!���YZ ����@��8A0,���4c�O�A�	���]u�,�N�Ztw3Ă<��co��XO7�j��1�?1�~rxR��o�=�APi�ӡ���eˌ��3�����	�ݎ�/�%s'ہw�x�ck�7V~��`�{��	��.؟���<��ی��/.�,T��0Rt}���;��Ϥ7ײAw�M��>}�[xt8s�ɟ��p�$5��#��q�{�ä����Dm�K(�v��q#D�!���x�nJ�]��R�H��;8��31�g	��W"�3��3�A�+��Ii�]T��=L����צ��5/�)�������x�G<���m�j��C<n:u���/��u,KF3�YN6��Z�ˎQq���nZn����㊤f���|Y�Z)A#�C�:��<{ڔ�:mr7F���e�»7G�*��eX���ס���O�T�4y~��/�z���nA  #9�f�9Z��p/�����Z�c����zҹG$˲b�f���jA���=�虫�H�����7��Z�u��x~�,�AB�ĥ�T�.;�ɲ3�*^H���g�N�h�Һ1�Б9�ֳ{�2��X����gFz���bg�����ea�'�G˪)�9����?�Z!���_�v������Kw�~w	mɯ�?�B����j��h���2*�Icw�ۓ�bWQ���K��Og�����Ӥ�zK �ʐ�B�2�J��Y��C{\t\:E���B�7�֋6�4֦` P����>����c�Of��Г%^��7�?,�.9��D�[��Y'�-z�\+�ḧ8!��u����㛣�Mh�A�\V\O��;kh����g�/"�_z��d@A6�C3���7��S֩��K�-DӘXO|���d�XÁF6��˃��t�t�`�4�ɯ ���j�ꆦ	�眱I��B����$^9�$Z�����¥#�z���K6�CY��@R5����۔��0u⅑��zO��K��-����S1j#ȸB�f�H;ђMe�2��&� U��#��� #���`~�Ȓ�R��1��*&�15s/��|���5 �ͥX��=N�8�}f�p����13���{P
Kj:�ćfl�q^ϓ8d�\ēޒWC��.��Nz07�d�d�~��tΣ����U�Z��o|mDШ� �p`��{��R �B��}��kN66���xXB���v�K�u�:7\~C�e�z8H�c���fA �.�Q#0�����
�Ce�
��nj�v����,5.H��@�����*��o���˾$H2N�����\��{>�HӮD��%@�u�,#��
����K��|B�6�A����^@�aƂ�ˎK�\����.C �>C��}�Bd5.6�9ad�H��wL?󿗳���[�#G�]��\T@ߑBC�y���A������7��J+��J�=_��/������ŵXn������+�Wb�ܻ��Ҟ��-��;�Y/+�n|e�t!�PR"fba��Q�~���W�
��^0s���ra;��
���I�I#4,��J&2慺������ב�i/��[\\^����m�A�XvP	���o�ѢZ��:���F�6R�^5��yn�gX��%���Uņ��C�FC���TcY\]��il25��Q��4cm���Z�nC�ݥ%d�iq�;���<�km��l�����G��Y��V��뼻���7<����������#�~������,·�?OiAu�7ۥ�{W�m�`w;2"����/\�?7���ƽ���4A@�~����2^��ueTT�����1;�^;Tv��5.�4܆�]�3Q�g	$�Lf$�+ ����"���%b�	��:����w��5�ה���;���%FЯkK�Q,w�&�`�t~�J��ﱛ�B�ltc�4���%�±�2���d�h9ֳ�B����l�����UG']Oqw,iv$ߝ����j}*�b�8����"�+",���\)�:�`f�qCb(�����/64+r/��u�A\�z�> �41:Pt.^o,�?"�*�Zh%s��5o�Z=�Xĺpm�D�Ϯ_���|1;ځ�H6���#��ݰG$
_M-��4�m̭���1z��H�X���c�X��W�t�v���~Ҷ��Hs#���@ri7��`��	�1��]p�Q�E*��q%��E�ŒDLb���ۄ� 6X�^����ϝ�[�ZR@j�%��pI�XD���A�g�:5�.;��$�n}c-�;6I~� �a�O��^[+����j��f�WE�	�o��#�zr���
{��PJǵ�;1���c�4UH�w��� ��*[�c�p��bI��p�"Z�-?���QgDa��s�.�!�a�唃����{Q-�_ՌdG����:��@+(���mo��,�/�pE6�t� 6hr���,Q���.�8i�kd�t���M6�7��^|�{Y޹<��4�l�J�����H����=�i���7��U�*T��[e��#�~�G���l'C��������d�41�cD
��E���s��h�d<����t���Z���w�eu�=W�^2P�k>��ۄ�M���BƂ,����5\�My��%�7Ѩ�3��(*��ђ�{@@Oð�X��.�Y�0�2���{`l���"�cl: �u��õz�����pD2M�z�hl�'��4b��pP��F�ع %M8�! �lA���?����D�×n���S��b�����Q�Þ��Ɉ��4�io�h=?Law�+/	U?ٽ�ןy�W�zl���#vr����R6sK��!r����_�ߢ������)
�����h:���UX��{��#,�_�sB;~�eGq=mʩ���SC�]���3Z�6���1����L���~���f����pP�5/�e��H�����MCٸc��x5��}F"�Ǌ[�2О�$���《7<N��]�B��S��������|��b;�:8`�jE�>�'��vz��ߗ�J�(!ih=��e{ե�቟3��tl������5�E�V�#1l�}���`�oIc�e\�����?��'��tl��6�'��NBX��5���mN���'��.�6`�7A��ړӤ����A4��Ϭ���Љ��혼�o�sĆ�Տ~5�-q?���`�1�D��^I���XҌ4�R�y�	N �wxgP-��"6�a��noX��k���_`X����X�`#4�~��%���8~'�n�q�@ҰL�4X�M{��F��u���Ng��T��rV7�Y1���]��v_[��Dz�`�g��],g�A� �����������,-���a1�4��}Xr���P�A�����1t�@J�fu�k��K��V4��w�f>>JX�Fk��КMh�gY�suW�.1�u��ѓ_�дˇ��C�9�i��C��WˎԾ?=>s;�p��pH2� �b/�Vn+��X���>(<��}c��s@J0��QC���E������{^�������щ�ey�A�#icn���ݯF�就+WO�Qߨr
�k��fm.�I/'PYc�On��i���F
�_E�,�ㆆP@l ���N���N���X,�=�	j�X�Z���:ix(s@8g��^��m��)�F�|l5��F�����-�AI�	������5Q"m���_F���Q�A4o��^��D�GG�1�BX�;��[(.����ep��).�n�N?��7���ڶt�PL���<:��$0$�6n4����=06��2�Y�z�)��Θ�|:��f��%�۶;�������'}����N�E�1���j�Pj����,�5���y;��M�/��e/�pF&���7QbH��'k�QSO����?�ߙJ3N���Q:�~�����M��^B���H�J1A���!�Q��>6};]<p���G�� ���쳕�Y�Z3�S8��r��C�bM8�6p����ӛ����ڶ�sd�t���|#�O����u~6M�M�8p�`f�l�Z����{�Y�tjF��ym���2��	����.�s����8��{�<������I�ȟ�x"G�ĶWF�/��yF�6p2X͝�ί|�aĦ�� �8�����9�W;8���DY��4T$�7�'�'���NcY�r��i6K�7���tA#�ii��;�Y�p�mf����&���%�N��*�������p�p��P�"���%��3��x��[���,|3(��&��%)a5_��
�+���30�X
�J���p�I�}��E�40��Rê?-�R8���������Kf��NP+�&�syzx��u�
g�{>��8���y)T���Ή'��`����\�'�⃝5������|αgéjh'�N_{����w��n8���ib8�0��w��J/8^�A������Q�ē�P�Em�?OrCi4��ZZYO���W6;�����|lLsߺ�8!(�D���uf8�3�>]_C�s�$Ґ�����3pb������������k�3-����Z�����3�F&�e8�f8�2��2<pBi �in��3��<g���v������x��3k4?�/�Y�sU8!��<�׿�'?p`ÎO����s�sK�=���;,�O8��bd�� pq1�`�F��b�3�n@�+oz�|t2ճ(2��'��lc����C`���n8�D�_��q���m�3�ez���1��ڐ������g��yP8!�p\<�/0\{�L�K�l.��cd|�F�3\��p2�p��Lp�fX>��<p���v[��ظ�a���C&8�<�P��6pv�Z]t9ù���PM�?M�sڒW��?B����X�|����o� �4n�m���� ײ��U5�;��u#s��N�?��Ͳ���� j(�2����,����j~y��%�8^��MSgp��v�wx/�����1�B�+i�/:_�{�	��=ӿ1�U	�h0�k�קѷY�Χ��2�����5��=��� �,6��(梭��e{�VO��ڨWD�H�L��W�v�#�n80ְ!�ŏ���x��s��pb���&�S0����3 �#��pl,��κ�'O#+��^�g�)�`8����`�8!+#��ŵz���cO�X3��f��/ȯe��ZR�N5Á$���XD��չ�u���'ng	*f�ls��<�A�pL�i?�7�
�653������W z���z��a[�Kn���hM�_���xw|1�fOˌȒ�@�3(�T�<�Z��C3W2�"XE��Ս�m�8��2���!�%"��>����nX�$p*�����@�i[�������`����f��o^�ڲf�M�	�GH\P=�w����#
���?�-���\B@zJ냂Bj'��Ia���� r����E|�H�,��b,Hq%��g��]~��|>��q)<#�����`�Yt�&8� n8�,-���d��L��p~b8�&82Q?���AL7�x��#�=����$31 ���_){`�p`���e�;���ہ�|:��q	<,�3��׆tgX\���h��3�y��,s�{���'���|/<�"��,��$>(A %��xW��7�����<���F�F�%���VoH���:�vXW�� g%{��Of7�'����.���h��{wguQ��q�)�7p��Ď�lbN��ء8k٣������	�*�F[p��d|�ء8�Kb���^t�n8�����lci��Ӹ��	����N�����( IS'�p{����6�ީ���b��v ��2��p$�鈋�7�8�tg9��|�t�u���Z���k���v����p�9���	���B5�?:�Hƻ����3�r�,��d��;�������_�/q1�x�<�%,�x �&�eq��3��sG�&8���DN':V��߯	�pz�� )��V0�s� gs��0��t�g)�s�-�t]�K"p 8}Lpv��8;��	�Z����ւ>.X��S<�XpT� 6�nD�����pY�{���y>��
�8�M��}]��a8V���8;X�|̰�
'��� Ə�[�lL�{���]�2���tr���|k\8��u!SW\b<ȁ!.��[�����/8༆��hOp@xS�Ϗa	)�=S>��ɲ����|���>NA�?�u�W�ko_@���E�p�'Dj
��@n���)��,��`��z    IEND�B`�PK   :Yd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   :Y�]��N � /   images/907530ff-a8af-4c9a-ad67-f4101e76dea0.png\�<���?�m7vk���Flڭf�e�!�]�m5���J%���ӧ�P�l��˖��\"�k%��E����0Hc�����������*3����y��9�׸q����/v~!$$��_�)BB�K�����l��t�5}�>��;-_A"�E��?��Ղ*$$������iS��7�g�M��{��y9	�h4ŋn.T�sN��^��xZ;���:���i�������`�RaGo������oޭ=&�����O��)�ʓc#ʓo4B���&�*��.���C�7l�|�돯��b�z����+��^��kY����зR�k�f��IB��>&"↼y�G1Y-nG�W�m����)����}CVܔ�������I�
;nX��r����K��}��	VYN#����� ���V/��)k���rG��]c6���h��S�T}�CV�)Ly����Z�li�Y_��ū��n^���LL�JH��t�3�h�=+gfR�g�n��k�^^*�0�K�����W2R.hɘ�,3�8�K_ZY�&_,cqO��mW�!'(2�:,I�1:嵆�����^��S��I�������[���^�]�Sq��K&��$M'�IVi-��ۧ��)Z�w��C���w��7����o���>��~�z<���h[[�aZ�z�7��0��.�6������AW�x�z+#U�v��\��ڵ�iܲlzk��Vobbb�J��������$jp��0v����K\Y�+7n��S�1�4{;��1�r̒{�Ai���o��z��U&��Kq�,�<O9�򱪴���Ɡ�x��_7A�������TU��s�k<Ե����)��Gs�)�p�l��U����_{1�58�
;�譓���y�>ۈ�j|�MjBB���i<j���Qe>,�6�h����dУ�mh��E�Q�����Uޕm�S�#Jb�U�����ըL���賫��2����O�h�M<b���%MtW>�njjڣ��#��	���.�A?/�P�o�(��(׻�����Ǡ����?��*����Kݣ4�4í��)����I߈��6�^#�߾}k��QW��X��4����H��9�FwN��~m�%7*i���4��e��5i�X���]_����G7v�L�����JP9T�1�s%���b��A:�k�\�HR�]J�~���X�,�<`n�]vG0��+놴�x~}��D7x8[<����=ޔ�D6�0�#�f�?;$����*]LMMYѻ4!�d����E�_�e��-lmul�	'H�
�7��F��}d�+4B��U>=���]�>�o]48�\kK�kva���zյt�7�&�0�!���ۢfôs�^����)]|zk������I�*�<L$K6��|w�מ���<��F�ݍ��()5��ώ̽�x����g�2�27���a&w��LG��a��N��p�ܪ:�Ru�)��Hw;\��I��%_��8���8�hڳb�A�>R���4w-**jϋ���S)��\�O����)T�3D=��#����d���t8�Ӝ*[�g�SZ_��������b����7��z�Z�o˾�/�gxv<��ܵ�^"99�����Ѻԃ�0!F��&�k�����m�K��{�L��߸��V�).ٹq�S�TaG�m.��͍��=���R!6�{-��%�f�Ҋp�tAs�%x�oZ�N�-��N2����ݻ`W�"~�������N��E%WV��N�$�D����ip\H��0-�����,u��/[f}�ڂ�[J�2�!A9e'�	&$mi�zK����p��Ǳ�3���B� ���r���F=%��ꐠ�����\=�������9x�o[ )���tE��Ǐ�,M���МL{�JǏo����Pg��f�'`��6�٤��mMH6ゥ89�Ǳ6)΅]����������{���x�<6@ou�s�����԰{��V������~�*ی+ X!��ge�?t�޽����.�i�� �{1_P���ޞ��s����.�?�z3"���7��,��# �6�GBh�1�,!��<�UU��7�����W'�+�5�4�q�$1�ꗖ�4c#���&K��s��<�
O����e�l�����G�·�?+��t)�a��FżO��31�2�w)�Gk[�?~~}J��)��\\\Ģ���1�I��!������)�忸e���1%M�ͫ��Y�M����������1�h�,���&h�����n!ebBweI����cF�dc�]��^k�x1���+I�F@ȓ]ߠ�,�*
����t��2^K�lPv����{R��a�K�� �T�R��&d�O�{噽��K�g����v�Byv�I��/)/���V�٥�nX
����������cY�`h�r�n-�\�WG�A�.:����� |]B�
�g�N��?�T;tHf��gM{b�}�hzir�����]>=b;v�8d%��r;O<�e��#�z�l��!q�v���N�S�Hq:��rp����<�����f:%�}���F��0myN��\H<%`䮹����,�~}ST��g�uu���Ϻ����,'s\����"_$1>����h��>ڻ��Ł�����I�"�Z��}>=򳳳qTf�al�O��K����
�qp��'�Ѳs��$TaZLe�Ҩ��)��Is+�يx:�Ǘ�{�Ոx�-�bk��{*2����&��4�dHb0���r��=�`(���D��ӧ���W��kݦ,���}"4WEi�%>Sy��u�e=���u��}i޻o_��2^fҬca�-w��}_�~F��<�g������gΜ������C�^�6)5�:	�K,I�H\?��������vN	B��e/�'�u~��dQ�}j�j�J����*���ڼ_.k��꾵��+m�-L������<v�`Ne�9;J)N���F/g�oP�ٰ�ߖ	��t�Ѩ�)�t@A�2�P)�0����ô�u[�A���K�?�m*�#�@�M�Ux��ͼU��;q����1�\[��B�@��Y��o\��H�؎���0��#Ii�K�g"G'�{��U=�h�Cv���PM7x�6u5.���ܹ
��,�� �\������4sብK.Y�Xx���%J����ĕĩy3����S�o�{1�c�u|�q/�<l���8���1Ӝ��c�#^=z��'�R��1i�e��<�]�%�9�"!t����Mp|g�6syL�e�\g�s���2iv3�JU�$�(��^7�:�����t:u�l6�Nh�z�<�$>��'�ϑ�*���u��ŋ�.�!1bj:�����r��;$$r�x�O��3�؏��c��|�)�������L1+��%�}���\�����1>�D��t����US�s�7�y�����*K}O�[�Y>* Aa6��4蚘������G�9So�`	�3�ʸUL���a��bN��ρcI��C�_ZO]]�m�c��m�mف`y/����s���q�#���y�����H#{H�}.ٕ�_�.� �����h�D �l1]�8''�F����n2r���Lz�A�������2��#��L�M�����;&!h�����$��$%##��o޼�B���%�_�h�c����2��O��>C/O��"[�I�� �@W���w��k��RJ�>S��K6���b����H��!6�=�>���������<��N�7D���LI���L�Q��?��",VRNXl>3��˅�esC���^k��p�MlX��h�D����
�Dl8Iג�𛾴{�d
*KM�*5؝XAA�UbU�u�R'�x�pa=�	*�zu:d$ɜB�KIM]sc�#��i����7"2����F�R���)z�y`;��K�w�
O\�<����Nu��""l�>�+qO�����Iԧn����0�|!'����
*�T�C-<���a��yDbLA(��j�c�J� 2�ܟ��ݟdbB�0��|����48���w�;l]�e��%/��������#�����?�q�R��g�-C��H�m��V= �������PmO����=Ω�����	}�ɐ{�&�%�qa����赹�P�!�R���˼G�{N
;/��<��Ď��am�a��]J�2�(��e��aB��^y�]ys�������h�KPQoG�X�K���]���1a/~��b5�� ��Z>����'� 0|q�S��ۉm(y�FM���8�������pI�mh�ak8_���$%-��f�\^�����o�UJ+*��H#�=�W�Nj���cr��$F���BE��$���܀�5���;��4H���'NOB	`NȂ���ƿ\�������XȌ��+��e�v�֧Gě�kC�L�z����`0J333���dr�m$I$�����ǚ�މ��p���W���� �ڊ�����g�ӓ�����R1��� c"���k}I#�uC3Ő��b@uf�ͻ�>;77���E��x�s��Z���Pc&k
�{H&�Я�nddęL��C�M�7.}�I��K�DTh^�,Uc��<��LK.U\�������,p��]�['o_z
oW�,[�5���~Jd��x���Q�m��<WK������&	�O�BY���ӳ����"¦W�䭴!���G&I�ۻ�����#��}����	�_;���bZ��bI�ʒ[DG�t{|z��qx���� f93�J[�P-�oK�i�{��俠ĹQ��w�`yaA�d_� �N)SVS+~K�඾�;hyR�*�U�M��d�#L��'��?� ��ԁdw7DU.��f2h60�nY�u��ݎ�jS��CU,�?2ݵXW]7N��~�5Ч]br�n~%a�{������PW��c'��KߒIJP�B�e�]8��XM����3�溱��lK�m�_�
Wۆ���M�� +B<�<a!~[��\02˧' �l�V/��nݺE#XgY󔽉��U�Sn��~m�nX2j�1>f�Bm���)"i]bv���%��֪:%ޟC�Ҕ[�[�[[�#JP���sRo�AE���{�B����G�/�fՉX�%V��fQi�B�U���0B1хqH��Q����b0����ej���- 12�I���jH�x���bJ`��nc���{~@�1��T�h�@��J�Zh�)jY�s(�Y͓��w���;jp��-�
Qtv�G[D[`%�7y�k�vuu�v�e2��ϑHM��d���qq����	LH5������.�q��"�~#n�@����'��}v������;d���P�X(.n�P)�}�E��TВ+�o�QUU^YS\���Gh��UN<x��x�[�������!��t�b��~�[I�����8`S�BLu�Dk�����BC��j�na�}�7�T��f����0$�Q�'���ږm�����!}�|HȪ&8��&���	.|���7u��3��1K���ŚJ�̯5B/��x��B��(�98�������1��R)P��c킔��ebl������Kv���B=쪟tu��@_pd58[�j[[ۚa6 ��d�Sb�é���
~��f�8%;����g|���ʙ����ՑU��	|E��snDTTU�ޞ�[���ñ�����RSSS��Sgb�����6�����4°���4$�pWG�	�./����T(���S��م:qI?!��'	���gϖy�C�����!9�V�I%�rg�!Y��:��^������`0�+���%w*�~�
�(Om$)\��^���q��@Pb	[z�]�Wo�o�u��Ԟ�4�NY��\}MESs��N/�C��
�V�eH��ܒYi'�(R<�l����N���I�;��}�a���;`�pb1��x1��qw�J�;Z��-48\�s1��~��?'6ӹ�Z查U1�U�'$��F�0L�����i���"�Ɗm�s�1���پ�n�p�C�/0��la�YR��I��^^�MR�J�xd�)�h�:Š��$�N�n�{��Io�RS���K'	�HYz��b���Vm��z�8�t|�d���\M�ޏ�׌�>�mM��s"� �ݤYy�|���*5od���]����I��v�Cm�1w	������imm�_�V^�cf=��W���g�b�Cs�K�)ZH���������Kh�}H�*�˛f��-������_�s����B��d� �<F9O	E'o���5Մj	4�	t�g��C�,�Ǉ������{�s��GbccG��ӫ$�g����^i�Pȡ��QP� r[ab8ͅ��v��%�.��	�	�8�A��$�� .�0;�	C���Y�[�_(uX�""�pN]m�'r�nc�MP�uזk�N��u9��j�y+�%;�,b�q��N�,�`��z����2a���$�=JEX��Wyt�Be��P3�e�&��÷۱��dKD��m��F(k������4�1�L�W4bQJ8d�v)ʥC��\�n�~jdj�P,��j�J"�^XeC-�H2�J�_��]���)Y���)U~l5oN��%x/0�X���@�Ν;v�Z�.�Udv�xJ�bmmmj����R'�W|��nag��&��-j���+�%s 2k��);�
v��?w�������~F����!�8jU"u� ��������{u{��gQ�G��L�MY\��Yh��Y(=�����z���g���G���7��$����%��y@�T��h�u��^�r8*�p�+G���*55A�?�)'-�Y�8�=�R�a�2IMZ���>��k����^��ӓ糭&���W�9��kam]х��$��ĠV�h���\�FaQ�����ur�X��1�CR��������I*6%�Y�=;�K �K��~������Eз49B��V����Ntr�x}�ZY>��/
s�eK�"yv#Iv����D�#:�ؙ# ��2�;�	�޼	�����X����b(Ƭ�\X���x�լ�hr�9�7oV*EH&<����ޞq)�:��>C��-i�FFF
���
��#��\��Q�����v��	�G­�j%��oxe0�0MMM���e/�+5�^�������v�e21���C� �,����nk��������]o݇N...1>6��~"H/5�[�cBFmג,�y�Z2}��x�sss�fD��H#S���T���������)��7�e��gI�^�F���)		��T��ߋ�X�C3hî�ҶQ-+��:_v@M�������atnoI}��J{�[9���2��(��룃���R/��*����[�(��#�����9ZƤ`lR�(�l"�,mw�X ��!��ۯ$Ƌp1]m�}nt�6V���([���$\q�]����ƈJ�O��3N�#��S��r�E,t�E����r�%���~gt����#�:�ʆ����+�eQ����
;�a��H�Z,�%;�j,�k� �����:H0�rEu��ƶ�d���+7��f�/�|������<�����b*�in^��*N�J�'QK��?��6]UzkI[lS� ��9�|H����h�9-�;Y�p��Z2�E��\�-�oj�Ֆa�[���DH�^\S�T9������߾}�"[�k���
q=�������~m	D��T�v�j��7	�.d�%P�@&;Y��9�dQ��4���I1�D�Rv!�ц�
���e��U[���Z��AQ{�-����!9�Kʒ˿d�`���,	��Ҝ+��%8���<�V���͒sx[�y?���_I+Ÿ����-n���l=@�sPSx��VBBBs%݊�v��� @��/��3l�4�FGG�b�s�(oǠ�����;.���$*���Oe�K�ٚ�Y����E��:;B��I����Ҋ�����&�P��B*?�9���\�ijrJJH�O�h+T������䖝�~VnO��CY��=50��!J��]������>ZZ�T���_�1�(�եEa�Ɏ_���H߃�X�Ш���0;���t^Z�Կ]�݌����N`�H
�tJ�O�1��-�΍ַ����TX���:3��+	yj�8��T֙3g��髦�o�Qd��R�F�gI��[�1�e���k��*~nRtb'��l�<��P�-6mK,����[�����+�4�dn�m�La�a-�SǫɹM9!X�I"���l.��R�����R����X����KLL��~E�֜�pӒ�>$-j>�.-�)n��(Qg��
ǹwj�����i0ߚ�~�i!�������T��q>Ѕ@hI.)��������� W�5��mC��!�M���19�M��N=�����ļ��WYYyXZT-��ʮ�n ���\�	J�i�a�8��l�Tm�r���$�����������#��-�֪�¾�f�l^mħ;X{��1�E��.{e��.+i~��*�zA��"�;ˍ�pPZTBe����ˠ?���3ɩ ����Ą�%\�֤�y0tY�1��cWV��'��<Im�4����:i@�C�f���A���a΄{"R����b��,����ו�ħ`mF��o������Es�X��Xfd�q~��+>%D���f�@��*�T8�.����4>�/ضm8~�U�S�!�]Ju.E1'c��Z�Z\|�����!��F&�
���TD<8~z���������)�m �����D��o���_�����me��|��ݞ�[$'�c��ܤ�&����`��1�]��ɈW\�Vx#�7���<Ls1���$K<{��s�ja֓��rqq���X�\�5�Kb�.�^��#/�/��K�8F�^s�>�i��O�4֩�ޚ\����i��*v]�ܝ��HR�Q��k]^^��<L��}���qP=�V�~�E�d�+�%�P�=�0֔�)d���b���t<���- [dEv_c`WH����(�t� �\X}��_�E�q�N��4���w�SL����33~�J][)��NE���lX����֧���ws����șM=�m�,�Z~6>>�0籌B�n�%K�9(aJ��+: �uO���}�.v��c����gϞ�D��܇y�s��RYի�&:��)Gͦ!�W����ڡC�)�ű�T��T�mT*՝��,��h�700��Q]�eFa��|V`e/�ZcQO���,5�rN�O����ڞ�D$��WVj���V�i{�$��*���V���2j�I��[�g�-zh$aj�q����q<�'��a���
�Q��e%6�<���Ȗ���ac�vP�40,�Bc����gmlV(<
чp6�����!/}�$93�<�����\�df)+X��m�d��z����n{�m0|.a��
����	�m�g�v�|�tg�u� �@���T�-�@V*u4w��΃M�41垬� �kӚ��]M�5-�҈5��$E���[NU{Ѷ�����!!�w����A��]���W�r��Bm�'�3f_/MU�y��Al�����z�sÛ��mE'n�{RR2_�Uom��KIZ��wh�k�!XNpC�e
ym�M�jh"v���EEs7�rt�;&�u����q�t�˯�h��⯬��:�61�!�u�0�ecQ�RDć
B�	i�����xGNW�����'�פ� �hZK�aZ��H�ކ�ZV�b���H%{7���O�qR����n*%�ڧ�(��k(S��<��:�1����b�9���a����D�P��7m��^�c[����[.|����������;�tO��}R���W��}4ͥ�1�y��6�e1�攕Y�v!#�vF>T�� �Э��Èև�{z�L��(����X�a��U[o7h��hT��9'6.n�j�B�����q�?8;F��}E�r8vm��v)�WǶ9J�������1"���kn�w�{N ���;����U�}�����*)����&�<��� ������mܵ���\<7�N�q��.\T�8C0�疭�H]��a���[XZ��D��ș��.,���3��U�!y�b,�� ,Z��@�;"RM��r���t��XFV�8���F��QJ��CK�ߤ���W�6�
]��&Da�	��)��
�Rh���`�u=wn��dc�e�ht���-�Pgw�)��*=�T��z���>�&�
�|��H�����A�O��]WBւ��Bh��21��}}k�m_�Uj~���!��ݻ}���į���.TS���d�|�/��n�)�T_t�̼��e��Z�&���� ��{e��>��W8��y�?:pq,C�֭[�
7۱yd����ҽ�|����n�i��P}T��0��ȹ�����<vi#aii�ҧ�tO���Z�@��������6�/�����I�
r�����|�{E�k+�TN���pyW��:3�rĭx���zy��	T�? ����L{��܅��s���#�Sx2���w?|�����!����bA�\.7f���3z��ҨOy���/�|�Cd XH	�rd�߻��o}n�Dh�B#f;���<�m�>v�+���1?�,�MO��ϘB����C�Â����B��@�쬬�r�GqAZ[P���5��^WW�w�T��g�����iYY/ٻ��^JB���n.r�rV?ڐ_q&v�=��ck��+q���8��!�ؑ��� e4�G �Hvҷ\V#��Ei�<�;^sS����0���E�*�9���"t�6�kwC�7�Pa*a��ɾ ��J�Ϳ �5sP���K�&����Z��_��T��x<]�Ffw���SPV�h�d��y�L��iTT�!]'��EE!D� �=|M�^�F�3�3Z2v�����E�.���k9�xc�E�6���@㇕��ǀ��رcGo�7s�f�7?"�t�^��2���Y��A����%��qZ�*oS�#��o=�İ�!�6�����5��÷>� |�CIpD��34���#�㦩Yv+��k�-�P6+)ˑ@Y�.�"t��k�YY!ܷ����yg1��_Q�����do���c��k@�r�����#��*�g�x����(��!��X ��I@v1T1��?�v�|Q�`
�,#�7��s�ң�Nw��`~��鉶�����&�V�D�Ξ��q$1���tQ��bs�2̞�#��8�Q�M����}s��7C?~�,�ɇ�v���{�$"e�I|l(A/�+H�5�0���H%*�����i�"Tpk�YпԓR�������y�*�qm�wC����V�/�~Wߔ�^�Dχl������+k��h�H3њ�=�Ն���;�m;�8��"vJIk�'B5O��>��r�F�����roo/+1��>vUVV�C��y(t1Ȕ�ТTb)?�X�>��/�1R���M����C�A��~�IU��N)U?��IU��0E��w�0-~�I;�G��Ht�����D	�ZM�X'UՂ|�@)ׯ_��\4���[c#���w��8zp�(�=�@���߭:��6bO���� ~L N�$x��o��u5��Xq��"�f�i�q�<ޕ>
���y)a�.��K��"(����܏+��uKE��nbj*�K�P�⵿�^Yٽ��j��R?
BaJ�根)y��n�m�		��;ru~��ч� q�d;�7�+p^sƞ
�����ɟhҪS�<��3Pc]�]��"H���,�����y�]l�0I]Mc�&�������2�6�5U%$$lC-Cg�h�>h�M]�r���]��"��W2��*�'��{����k��S�f��>������#����q����%��&P������v��j�q�m8���t��A6�1	�ȣ$0�k� � uL�QKR4�OZ4<�����O���)An)��Wq!�璣�P�J]��%�v�g��~f��@'�Ҏm֚���]�Z��%$�3:}roȗAm���oP�L�H~S��*��ATUBowHMM�=A!��
�sI��&6=tש�v��}g����՘�w�^�g
Y7���ɢ*����Sw�c_JA!����!RJ��5��prhp_�����Ss�;T�ަ|a�c��P�ڇ���8Ek!g�s=���n�X��\Yi�� aC��+��K��3vX�x�����@b %�C㇟p(�9��v�5�0��i	Is�c�5(ot<��f6a֪ǧ5t,{PalL�&�c	RTHu��k%M�6�&&�To�,��W��v�[*&�hy�)��C������)���>6		��h���C�)��� �AB?g�J��[�#G�����Կ�&s�$M�Ѣs@�U�]���g�ቶ�J<^H!	�ͻ��Z�!/g`_I�����[`��y�&7�n<��)z��e=���5szgL}3$���-��׷�X����	�u@�'n);LL
]�\Nm��4�y�N�D�"Ӏq���5x\tZ��V��@u�N�"���o�w�����]4�K�_�C�n�~�$��C��G��w�{0M聺��N�V�>�
FH]�����G��U��@L�A�22��*�e��a߼y��ٳ~O�X�S�^#�TTI;�k�!��@�¬,�7�q�Q����.AR���Q�75��--�2}h�3�Ɏj��prC����N��	;���^j5������j=8�Ϛ�+���`�PȊ�?EG2x{;�9J��+9i;(���7D?*�1QRP�Ґ�"�C�5�k�C�r�K����u�OB�)�N�������3I��Ê�X�W�oA��j��*5�a�����D&9��g@M�����V�1>��¿�zHu�,/��/y�u	e�I0fL����M5�˗�����=��_�e([YY�^Nݳޠ
e`
���Ƽ@�f�����W�˚�N�A!��j#P[ͧ��������`	�8@�8���|f?=O�ޕ!������&1=Oe�?�YsI��%����C3�_򔯌��T�,
�k/b����Rg�v��r�Ip�;x��*�pr;��\����I�M ��GyB!y�s&y�U����V�%?U�I��;��3�E<	�nnUL<�&�:�R�0ٜ.28p�E\�/;Hs70�pfF
�G���/���=��ZM����J�M���};%���\�s�v���\y�������;(c���7�w���*$��>�����֢�[0�=S���8�����2�TtJJK���=�i�W��W���F����!)����%��峸�O��L��MLZM�N��(�_7|O�F�n.6+�W���4�L&�I���N��͢X����"�,ɪy�{J�E��Qlc�R����d1ؾ-� !�c�@mZBI�\�m�f���7�G��Nه�Y5��@�!L�{r�K%��ǮVi���- j�	���%�Q�
A��D��ֈ�
;��%1T�tM*m78���(��߻ F�3~At͍%_:Y�4�������^pi`I�JU��Ϻ$��_(i<t��6�哑-���a>h�zI�M�87+k|ѽ���'�<�/�+I��'3�M�p8�I�ڑ/P# }�����)�(��(D;jkP��pc۾ޟTU�7�UZ^�%��0��}�3|=\��`��i�9�Zt|��-쁈̬K��7h[ ���
jN��&��)٭�$�~�F0�'���5��}ȐI�f/P�V���q��D�� �<g����)�,_������w�
�9H����E�?!4DgI�Ez&�4��,��l��ٲIBo��/=_A���s�:�wcT�)f����o�E����Z�:���;h���D�����KlYN 8b�qR����WHc�����J��98Db#�V�}q�F����w�%�K���<j+=K� �<�k��f����(���h�{�#�VU]	Y�Bұ"++���q��d_~U�ڵt α�c�SmЧ��| ��e���9��P��Z��W�2=���*��DaE;���$�����h���H����j%��~6&|y�]�܁ۚF�[�$�lCW����*��&�-�\���K�,W�	Έ�ה�� �ݲ�?�&����ҴKQ����G�+��{���#��XuL�N�z֖V��xIk�p8���;�G�� �B��5��N-��J�6>6Jü+i���S�yh#h����l!
+>��(Ƞ�z���(l�bfFss����_�w�ٙC�`!p�&X
��ZsS�����աV�F�)���茏��)�K�8i���[b�T1�\��vY%�tS�MW7�Z3Y���t�:�φ��Aho����UMi��k�؀�~��������
֭��]G�R�A�p��V�N�S�?�����e��\ mŻ�}u%��]�͐��KAy
촘���X�������R)�h�����Wz �z�6�G$B��ԐFe?�S���</�UrR�$�C��kL�o�%N]ۺ	A�q�?��?/tuy��vH������t8����=�k%����]]ށ����xf�yt�d������'}M���P��'�:kɬ�@iʚ:-!T��)�`)d�Ql�k�H�̋�+��N�g������	V���3�	%l�=���99�W�>73��#���:;�|�9���|a�P�T��)��)HD��:��0GƹMI$A���5*�v�8�<RWW'lJv��i�íz-\>S���#����^~}���2����?�9���Y9�����O]�8{�s��=���Ͼ���F_��"���-��P��ySS�M����b�w�=�(ľ��� MX����Ɗ��1�a4���G�L��*�q<Nqś<�`x���~�ώܺuk*��XU�\P6;;�{
�**Ts��`���=׷�O�w����ѷ?��&�/�.C�[5�����ZY���z����B��J۩ۃ2�ON�*���Uz������Ûw_������!?�u��6�:���7c��"�s?���+onk��{܁���ʏ� ?^S.a�V�p��8ӕ��`�?�*G#���I�Ckk��x�-am��QT{� ���;a���+�'ږ+%�D���q�c���G��Ro�/MOLL\*�wOݦ\2%w�����@�V��B$��X�J�S�������N{����/�|0�x^�մvC�c�;dVxٓ�m��T�oKB5�yb��
m���PWE�?���������U�G���R��G��08���<��Y� 1�SPP�dZ���V��l����z"�&(�P��:x���prr������Mrn�������(=&@&��:*kB�'�ee@��l���e^��w���ڲ)&�i,RX��i��d`f��Y0H=�oG�y��Գvv��< ��}0�c��`��#�SF�~_�J�L9�^8VV�"��@�柠6ɉ�-�E=�1�
��O ����R�7��Z�=���H�������>�bWW�΃'f�$����'�̴�j��uh��]}}k]��GT]o%r?>!A�ݤos�O��k'G�>I7�.R�����<����d�v�i��.��cj6��$�gɤ&e�/���o�x905�F���.//���:j��8S��[{���R��@R����b���U�;]Gܮ\ܮw�H���ǋ�H�޼��t#]�7�Y��.BG�Ð�Н�񄄄�N|���\�n��&c������m.�
^�07k����<��|���-��[*�#׆|i`��
����q������4�9���n������埽��T�
�r�5eؒ�^_��P�kw4b��o!��ÖtA����J?�v����Qv������+q�LR*n#�wc���R?�@�T`�Wg�������	oF�PN��l�?R�p��xY՚H�=Q����၁�&�	n��}׵�E�FMTs.t�=��C���ev�B�����.�00��;���' ��KNN΅�I���f~@�*l�Z�:�-u��T�q
=@�lto���:5���;&�0m�l'@�	�md``��� �����������SS����k��j��N�Nnb	�ae��E��a�L&��E��g��1>~LPu)V8�(���i`�9��e~~�1r2��2���R�2ۆ/���m���������Y 6�q�2���������h�()(�}Y�j�J�;-�C������p��~�e�*풖^�#9�-m��κ�|[	������:j�{zV�f�*�K?c�*�P�
��D���N���x��N�f�هYY�ֶ��wp�S7s�oٹ�S����7�`�[3�d��"���˥ۗ���6v3�a]�ͥ尸�J7��_T!p���Wx�S���/���߃��A� ߴ�~�~���Ļ�ꎢ�R��J֤/n.n�S�5>��x������)���%6N�T�5��׷>������[���v�Z����~:43_,���7���\�gc{���\���l�zc޼yc��x�L�`ȅFH!b��A&�z��-���:<I��O( i�f�&�ʮ�+�������8�7^@E�3j]:F��,)�\�w/++����L
��g�RySSv��Gp{)��>�M�n���ra����g�Th��z�����p�2��'vs��Q���( ��]
�4��@�K`T&��,=�/,�q�̬=!9Y�o�[f��^!�Z�!��D�P��"�9�e@0ʨ#��8;[�����q�.Ģ�x���r��ZIC�w(�`T\Tp L@�_�e�;������,��RS�A=%x4��6�� ��UGG��7z��Ϋ!7����(r�^��Η���従$j���@5a�s���89��%�VE���u]vϵ�v���o���������m*|�|��@
%�\��ɹ�s����֖�I��#���ۏ�
E�2�( Mo�;����{�֢ٓI��ɹ��	ߴ�]HLc��kT#H��_��X,j����pQ=�h�:^j}s�c>�����%q�e<P��!�Nm7C�*���7�M��ǎ���-�F���Hz����O�|X��i����?�]X��%Ĉ/!�B�{��D��f�Ft�G]Zt-����o��)4�(()A�|��Ԝ&���*U`r�]'����Ꜷ�y�F��/����(L�gtT���\��o�yxU3~A�Bc�����	����^��Ǘ���=��*�i���7o�PB�k��zY������5%�O���UmcZ��ޏ�9���8cTe�+�~m0#��ѣ%X��N�a+++wu��K�����)A�\@e���nZ�g���B)5��f��[6�9f+4*�$E,������V�����6�h�]��\2��G
�e7� ��}���\ݓ�_����=�b�*A�u�\�Ţ�����k��İc'c�����d�y�^���#=K�˗�����de�z��/�qP--�ǿd�k���?����f�Y ;�o]�n� ^C�S�.�3�����s����z��]�N��qMt`��� 1x����7TRz>a���ru_�⎛O!�\o�����B����h΃D/w�o��l����`*x78�>�"6���f�(���/�.�^[rfHӳ�3#	��
�X�B�hgX>��*SXz�|x	d�q��ͭzj41���B��zIS �A'�"ץ�M�%&�T���1�d��(v(�#���>�*��E+�r[�REH�q*wʅK��bb�n��*����c��:ǼW{�{z���jf컗�o��grK�8�# �ͺl퀡���_�I|"���̬	U�Ƭ��H�r톲r"(]��[qC\�&���_ x�s��t���h�Bd��P��8'�Nz�P�=��|U�B��om��U����^xx|W+:1U6��-�S>ഏ��>�A���N0�mT�K_���f�[mM�~ff�J�J~������*҄�j��P���ļ�����I"j=�HK[7��d���C}-��_��!ȮBR� ���1�� X��^���� `a �o��P�����FC�a�vY�T# �h�Glնa�'w����^"�Qӂ�tё08��×M�3G!aGBJ�Ȏ��ǔTz����GxrK<�Njj�������ȹ��?�V�ppq��㩂�Dw�+�>���'O�m�Y"���҅��C.�8��ff�P��PUUUj�y�,�Ȯ��s�*rE�d���7��������R��Ӳ����e��^�S㜛S�M���������5ϟ��L:�4o�1��&ж�(�鍉�8	���� ���ҽ�!?`�~�ay||ܝ�Z����r�G�e���vF����w�������_��p��Ѫ�,�}���v��[���ŋ���}�Q�
7D�?X�cf�X��K��J	m?
	}[���n=��u_�+��;���6�@Iǅ������-��x������@� ��9�Bd�r:��]�t\���u�e3�5���������7�ͺ�,~0 U$���TH� �{.�����;t�R�Yx��Eitr�����ߡ|������5�l��CzCV���h�;r�w_d�T\��Dڶ��ۨ@��Iuu�X]�Ԛ+�S�Uh�<��G�>�g�V��!҉<6��n|��h�Ľ��
Zp��n����}\ZQ�w*�P7�����\+���$a��,�s6�Kyk�q��
@�������_V������ˌ$�R ��)���kHj�$�+���q�d���پMW�9"���	ʟ���ǵ���E���J� q�+�~�X*�<B��s���^�M��gi��j 9�������҈*��oD!jxLd7�h�}8�|ޞd�G�(yo��9�l�ٸ$ݫ|���!1Й��I_	`�ūX�"�T�hZ�]t�fx��#�K�������`��U*�ME��>,R���aP�Q� s�Z�Al�P!H#5����j�*��!�"F�L"2÷�	������[�������޿��sεo���,w?H9/^�a8��x�fm��}�.��J��ߧ�5�d�ڷUy�Ⱥ�0�ځ��.v򣣣�٢`cĈ��]����{��N�/˃���+����N]�w�;�
e2�۱]II)B�v"�d���Wɴ���E�y��JX�x~�2��n40$�J?Ȣ��&>W�xl6���,K������_�$&%��W�4������8{�t���@���ym۽���/?)
��럵��T�_�<�d2�@�ħ�*M,��h�q�̈'�>ߒ�-�p�&lK��폸�I !���2/�u���V��S�����_�ۮ�V\R2o�TpP\^�����A�?�ltp�־���zW]&�@rE������D<��8��6-�%O ��0����[����By��@�<��s� �Ո�L)�Π�����|ЙA��	y���`�Y�-�_�<��7>��x��7�h<X>��I��e�2*�v��V��Jv>:�序P|��ˣ�.����M
�\&�UB'U~��oT�/[�tϓ.�C����|��T��`�����y{���B��h�'�N��\�f��ۢ)���]4F���]�qv�;�Ν1؛ׯT�0<��K�7���R8y�+$�uO�����腚���jY��@��]A5g��@�UcZ=�ؙjd��hxm�� ��W?R���I�0�S�5���F~�}�*_Yf��L���W�����>�F������+V�)�%��Krf��.~���#y}��N�:�E�K�X!�o��Hkܼ�z�Fғ��߄�9���>��zwlӹ/lW l�N�a0<�xh�f5�}L1;xkY��<NFG�t�Z����s��}���w��M�0�f�ɜ�0�8O.Ȼ�y���������ߘ�xϺ��孻FFF����|�2�`�)�`��[�PϜǕ�9�Kw�Mb=�GQ�G�1���*�TN��I�rURa�щ�gt���ڪؑ�)xz����[YU5¤�]��O��W>Ag�I��~�.�����2A�I����<00 (d�k�dP �9�*N�:���$`�C�Z%o Amu4k�VU����ŀ�3ʽ�_k�<��bY��GGL�g�]���Vw**f���X�Ó�'>��֦����7@0�D)��>���ZXX�j�ÆWY�]h�x5�>=;���AǺ+;cG>5���E\��a���w�Qr�p��\�s�u��ѵ�ׇ��U!��c�Ox� -;��6�~��;��+���o޼�?>>>�����rӉ6&�\�J�p�8�;-�Ǎ��/�1`�@�x��&�_]�w�ch�����(�oQSS�z?����c�[o�2ue�� �z � 4*�Z���t?�|�qoPಟ �[��IXw��;��܃�S�����ܪ3T��7N��i��k�6e�U���H�5��� {(��\>��bW�.��hO�U:+8��\2���9�n�PWIee�Y�Թ�Nw^�����@X��lu���t�p#�!�2�����(��ȿk�J�����9�$)�[����p/I��c��ٹB��H������79��x��&$��Y����]�qv�xOϰM$�GK�����o�r��n��R˄/�T�u�(���Rxl��]P�dY�z4�MHѮ�4y��	��+5�e9U��:���{Co���$����B�C6�%<��s�஧���˧zF&���$(lɘ�ק@_2���#�;�-qT�F<�+u��5c���!,�W\�~���I�:m' �/{��$f���F`�@���O��mc�����)3!n�:[0w=C~3�j����Y]Z��3�
z��ձ�����.<�������w@���-Yz�{��`�kcB	�� �T�Hk��Z������2�������O"��C@k���ܔ���sލȧ��0f���y��j��T�����5�k�u,�1}�SQ��f1D$uǾ�� Cm_����HNNNy7�J��D�%ݥ�?{���
��� ���Ay]�^����3���r�P��V);w4��ݒ��.��p�Pk{�UYVZzV�݃,o4�=�j XiL��H�m�B��׺�~}�FkFo��Z�Ж�	�?�S�5���'���wSw��ͭtX�9%��l\�ٛ��"+g6�O����2Q��
�~*\a�I'�5"�d������O��U�����)`l�/�+��8ŞT���Z�́	�?N���A�~�R��
Pvっ����q��y�}�?�R"GEA8��C�C-q����.������ʈ,|�NO%xɻ��p5�k�Ÿ]��+���Ԛ
��q�#Ną��8��J��p�N��^�y+2픡�Ri��S�CxO���c $
ۘ�i�7�Y;q\���yFS3�WE�.pK&/���:��^�,�\��lܮs?fu��� �Ԉ�\&�B1��^��a�0^:���;;�8Ac���0U�z�j	`,�m'�W0u&0� W6X�
b�K�������
��'�$�nm`I����W��U�P ��˄��0],	��K����ޥYd:�5
S�^+�W��H���]<��:���S��x��F�����r�Z��p.�Ķ� ��ȈQ�צ��n����B�{�6�����X�@�3 yR���Kf��XIWxCW��" ��NHagO���P�E\n20�%.w��Q �=ť�� ֑iހ�22�j�A��(�K4��^O)��w8��][Z�w��5K�������^�+Q9y�'���������!d4k�j>b�!688���N��;��.ƣ��ʀ��]�z�,ʉ'�v��7Y}tg��~�3k43�q��F1�m��<�D�R�&_ʊ�Z؎/�X@��܌�|�;�`�U�N~#̮D6l�y_����
: x��g����E�k�/��ѫ� �i#IJ�g�t���Q-�|4����ҝݴŬ��,��lL!lT'�;:f� ��A%�6&�G-/��];�G �l��LCD
		麨����S�W����8�pX^��/��H�Ed��{�A��������k;��	�Jգ��Kh����Z�3j�
)�@����a)�(�\0��\�氞m�S�6�3���q�r�A*����.�r�q��D�&�� ҄�i2���O�,/lo9(o���<���+�#�D�� p��<`�+w�}r5�eq�S:�<�*��l|� ��o���Q<d��T������������{���"<�j�/o6RĲ$�V�i������V��h���`��9i�	�fKQ���Ƨ��2���077'��[�w��;�K�hV��

�����`��q�5}�y�v&�LfB�>����{Y��mɺC�b��2�����m@�E�{��u|�/c��4@�ં�'3-Y6�5��*(�8 W3 -O\��Z���	4]<;z��g��BI|�m�B ��r�3�o+���Hmm� �fڟ��5N#p󼩗J
��	
�1����|��?�����v8�P��*��{[�@(��8T����A|�M�������@	/"�ޘ{�BK��2}%1%���?��Ɍߕ!����F���y9>�
ɓ$������-,�� ��N�-����K�Z�!�p4�OEiH?{hq���
s�3X��Z�F�9�6;;� U��9~؂�a�3J��o�*��ۺ��b����0M�z�e��5P�m�I�œ,(�Ҳ�(�m�g�z�j��!�bV.`0<��rI�)���\T8)��
R�Ѹ;%���x3 g�x�r_��o埫�Í94�Q*���:�4�*���p�zO�);�zf�s�<�d���8�s���pxA�Oim���徂!��f�d3���Q	�?�w�f����Ə(� �/j��ʠc�!����K�/��3��^����s&����{+Wd ��̌��r&��gg�=����Mۇ�5�������@bo�ڷhhi+�.�(W�n�8w���� ��}f6�P����v�o��i	0����	��h��>�w��QJC�Q�- S�L}F�ȨQ�4N�gQA'W����|��ԽU�DeI�N�1������0DC�^0r�������I������g�52Q�mdʰ:�g� {mp�̒l�rS�m��e0��ٷ����l�j����7��w�ꉋ1HKXn��F&M�+�w��)�ş|���W}��ƺ���=�ɝ�T)��ow���X��|�s?/�A\�W5���� 1`���`�w�8t�a���RuO/?�u�4��׬���.Աpu���x���'ʐF3;lR���ɷ�~�m�����#���% l��7��:^wl߃��`dq�4��������r5�ߙ��F@��$�8����[%u� �O�M��r�U�#з�?7\�/�ٛ&Ä�B���J�8�lfY���١;8o�ܦP��?ّ X��fZ�2-�Z��C�S23h�����Zd�yǽbO!d�NZcԗut~�u�\��*v��f���,�ikM��JY�zi�U+p��O��1h�j�@����t� ��-"�=��8��e�����`�[�=
�%%&Wȍ��o)�`E������p�F�k�����������澒�bD�6]���4W��;*G�vBD�l,ٛe��/ٗ�����	Q��J��R�@�f劎@b5c���@7g ���U���uZ�2��2G��Z���ۋ�gkCr�&x�ůpD�S���*�eP�{�;�i�R��N�8����39�� 6w��T[�X�<���h@t�U�-D�6��ig����� cm��[��h%�Y�����PU`PЄ�e9(g�`ߥ��:(S�y��U�nԦ��]%��˛X�i�����սC�����:�U#�2�j����L=�oMߨ涁�!ո]Ȥ���	�P�W��+��o,7�ڐ�M����UtU��`��%n˸ZŔ�X����+%��Cr��@+�+.�'����ٙJ�G�����
=��uK^�f��]m�֝dXi��1���o�L�k��ɿ� �b�o�B�}T�}�:T͞7cmUW,�8P�e�� �5�kL���R=:]}�¯#S7���=��3��kS�l�y_ ��� � �RM�@��d��$@�VU��i��,Q���8cy�wo�$xI`�n��AFe���F�"������k�_�㌙�]i_s���V�;��B�}���O@���������f��{|���#�����K��@dzP�eP��A��WY�� ��5M��HW�뿧�D� S5.8�{�|�/,�Gv��FL������s�$��.��Oච��˨�im|L��O��6S9�elA"�]曃c�8����u��8[����X��k[�q�@@h�\&c�9��T�d�.��OJ�.�5(G����\��Ayǳ`rpa
X����񨑾�6�(�ց�4�䷟�Lf�o�Kt�M-U�9�?��ywЦJ��B�W���ȭ)��n,��o��;��a�jJ��������]e�J��N�?�a:������0Nõ[��iH'q�����R�%�2d�6����L&D��ލ�.�ut6q>^ؓ�EO"�#˛�V�e�����,��8��3��L��o�3�޽{�����͠�KQ�X�1�X�t�����?����S�G���T1�/e��u�-a(k�[5����nH&o�5kB7���L�,�ލ+�B�?:��zyz���&���b�>��>����
 Vv�r��*�����cu�rn6�7��R��N���������8���>+�)1^���3������R�,N��df���X�{�R��hз%8?��k�;qa&(O���@ؕɖ��p_�K���ˠ�e��'��!�.P� ���U_�-�����TdzB��.�I���d�ŀC�R���@x%���k���M����N89�U�iD��C�X�s۰��X"��@�pޠ�����v)dq}�~�X3Z4�f?����������EZ�W�[�ٷU���=(�{]��Ş
tn��101A:��t1ʍ��7.��):Gܱ��\�^d�	0S�=��^�&�9���[�Vp�\ɸ$�P�mg�p�^X�<ܣ+v H�J��rGg=�����Iw���2�z�����K���n���ۮ]�N�?_�]U��Ot�SY�]�d�C�������@�q���������Z6���<t�'�����T�8բN���,(U����O��@`r�Qx��<\(˕.���B�[nL�$�Ȉ,�MY�)_�mh�P���x@�8��dq)o�ӛx��4y?`|0��|�#�=Y\�~���ӛ��)�M��/풦1v�1�˕��t���]��1�䷒DD(Q9��U-�Z����r7��FU8�2bG�4]0���0�W�}��wO>A�gZ�P^�!�L��ч�3p���z��9vz�ja�Xb�,?PJ
+3um�F�bT�G��>�����%r��� �پ�Rqy�t�fm�ї��	���咹6��%`���1m;�-E�M�ݎ��<�h�x*�݄���b�J�H���3���=��%���zkd� �!�ʤv��=�q2�z_�%��UŌ�Jl��s�kI�tS���b|]<�M�~Z���k�!�ם?	:p����U8ܩ'W77�B�q봣Tq�eb<������,��T#�P�>�|��B�,y��%��?BD�A�׃�,:�W��-琐ܔ��iz��C����O���(���t Um�R C�S��	�3��,�_Z���t`�{���2�/^%!�2��U��j0��������,l��s�~j�R�qQQQ�(ϻ��w�C��s,Z��C�Cn�o�t6�	��K��`׊�����SG����}�s6�&hGr�� ]ɽ/�E�F��%0�� �D>���4#�E�;����8ם>Y2GF�b�����S�*,�w�u�mh�i�4"p�����@O�h���%���Ρ �1Z��[Y���Rh" A/iނ��X�0<��w+�2S���;�.?��wp�����-����@:�w>�����N�j��8�sN�g7��*���D�w�f�&3ە��ϖt�]"x�m����nC�}������l�|�WI9���,,��]�_;{��E���`��t���Q����P�<B"K===�k�́H!�/�(���.>Y}�Ӄgqu�N���:�e�y���7t �=��S/4
��ɏ��݆�W�ooJ�TV�� ���7H�q|���д�g;�`�A߆A��pBLg6��g�Yk E�@�SH6>��q��r6B�;��#(�{�\�KȚ��8=����A	��AH�@����qi��9u1�lrP��<AU���[�S �Mf�nk� ��Ni�~��K��?�߽y:a
]s��MV�d��$r�O'Iz��t���M�
�V���$J��lc�]<����5 ����?	϶ѥ���Ubo3.7~JzN\� d_�S5�b3N�/�� ��O��&|�Ɩ_<ZQQ�-�oA�g����᪢��|�FEH���R\��F�l��� �,G���p�# 7
������@���3�/q~�,�w����tj�q��_	�����괞�'B�7�9��Q �e�O��D;��\�1�	�T�C��r��m��E(9*U  �	>1�KF��d�@c���
�=faȷ�{f�]�0222.##s�&������$�IBI>*�R �U7YOrrrpi���� �q�;��B�9&�r~�LZ}��;#w�R]�w���u�L�?ԅs,�V���j������Y�^	J$�7+�	IF��=�ܝ��a��P�q6Ó?����J\��M�kp�%����ʸ����N�j&*���>�;/����a*�ol;?�a=�*�(��C%��o�wvιj֞�΀��	��=48vǖ���~T��Ķ�d����Z��>��Z��'?���/Nz�[�_6g��<+T%�s���h�p*��ȚX�sS��z��{�<���������w�w���ocj�J<�22:����︿�|~Dh�L��D��:Ď�Q���ju=�w- ��� :=H���c݇Ǧg��d֗�� ����:ئ.Z�CY ������9e��Ci���h��w=˓,_��7�{h�1�^7X�+R���-��?-a�6�TG?�Q:ՈɆ�������� ��d� фd��Չ�*w0�O�=�z�v�pt���gȯ�Km���U(;q2�����pk����W�;.h ��%����ꁣ�hu�����%�?�
���C3�DљNU�άt��-�e�gJ�2�?R�n�G������cg{�Z�bB@=�< h/��I���W��s�?�Ǘ�>�/���tu'Z���=YѺ�{5g'N|�q����8nI�d*eG���@�_�Qe���0O�����%@�p!�0厫j�2�!�v�w�_
��ne����fm3���fm����v�͘ni&#�,$M���m��I��)DK8��T�eԬ�
/�ؓ�a���De�8���u܍S�)���l u��y��N7ʒ��~JF	᭓d��Pۘ�96<�g����{i7D����x�2�D��j�S�rT1j��o�� �@�_,��i�i EdE?}��_-�ޠ�4)k=�)~�V��H���#��g�k�?	�1]|�U��~*��2k�~Q�M�]��г6���m�|���d(�,g��o���F�s=c㹣�ć|���͆����������o	-L�-��&�����ޝ�N�>�#�j���/i��u�����ݽ�\�;t���*��'�"IJ�����櫛m��b���?Nφ��%�*h1�U��b�����z���@͓֙{�:7W��w�E�H��O̗ũ�2�^e r5@���4|ZIy���|�rʕ�YLd���ލi_�;QmsJ?5����Î+�=��D�؎ѲkP���k�����3�i�.�ZE�(	ᓪ��!W�>y���{������ �>�	���H`g�S��ե(��sVo�ݾ�ŠJg�$@t<	S��vJ��G�Oij�/��Um�/ ���|1�U����u��g�S����o{7j<c�xͽ���e�L	��,D�.�D�y�p_����d��=Mޠ�೎��V�N��U�^4�P���rgձ���3Փ��^*-�*�!ֈg|}}9���N��s�G z���K���Āv�Ş�R~d�
����7s�C&dI�+�6B�� q�1�A�P�1P�}��V�]��b#]=��_ɳ���7LܱՁ&_�X�i��p� @����T���ů��Θ�<i7m��2-ŵ.��}�o)���������P�!�q'�3&��'��=(�/�RS��!Y���'MxJ3��}is�y�S
15&U�s��1��W������ų��^�-^'�s��~�0�Ŋ=���g��Ņ������x(Z�Oe��A1�{��eJ�h�;?�6.�'o$u=����!�?P���y�T�vtR6��oHk�yc�cPu����38sAO�=������-�}x�V'٬��ص�ؼ��-V��'0H5�Vi��咑�������y�u�6��\������Ş���'a|��58r~%��{���av�ǜ�)�.D�u�>ٜ�~ك>���F��L�5�6�������VVQ�$���V��sظ�����#�=�ʂu��gPpt)�-$uWR9��%%�ѯɔ`�]ŵ�^_з+����U0U��ԃ��[G�V:��׷Lp6Ğ��W������_z2+�,"ˌ�y�Z���U\@�| >�h2^��Y=���2g���;��k?�0���KU4��m�֝��]S	8��s|P2��;�!h���j�J:񋣠�*"��4�­x��g�X���ԩF Ow�s�2(�OQy��϶i5`�=����[��$&�Y�J��xo��ܐP�+5����/�7N�q�-m���
h�1�yC�B�| �b��kQ��+�r����ut���N5cH��+�g�ݻw����Z��a�	��ac�J�~�m�	t8y��3�(�����V;"o�fo;Y�L�`�J~;���[}�/_�\l���ř���À?~��Bօw�r��+���#K�,�W�ݻ0ݾ?(�]9����K�ζ��T�
, ��c��*��U��OS�+�FA�e�Vra���D��}��]1bV�x�`rj�T����L	���-��/?*���P.8�����u���Б�Y���ok1�'M�W�� 7�0
C�*(�8����7V��$�ʡJ�hr�X.����2}�eyy��G���r�e���1�6p~S}�@Oo�`	?��-9*��p}&�/c��N�@s���uO��X���4���1�s���}��$�(�/���2��Y���n*���{_P�_~��PP1�mf6B�y/�s�ؓ	�U�9~����'��ekJ�=����P�(�͏<e+y
8c+��R�nC������������L�_����|/��C�;��C�`�N
{���Ϻk�T4I��Rp��ڮL��X���"�Z�[Z[[M�P�$�,� �4������e�O	���)�V�C㝪�� ���wh��2��'ෆ;�,�Ğ|X���	�Ne��l?MN��~:`�R@s�բ��w}I�dsX����
��$����%C��JFMM-r��rS�'\o{F5H�Sr}S�k�����y�~W�ůs�� tl�>?w�
	���6(�~���Q^���!9�-r�W��3�޺����ҶJ+Fr-��%�����zÍ�D}��bG���Y��Ќ|b���MB@�#������o?V����nB�����,����ۗ�<�+ w�at[�Z���#	�����"���H�q�&S�m´
�B�{$�ᤷʚ53P�v��K�Ge�%AF�v�a[J�q�e?`����N����5��r��O��=���}Ͼu���H_|f�C/,�6<�\���F����Ľ�#�0��,d5(EhE
��7`�8 �5����I��m;��Rt�)�A�^�'�QL��%jTM�g�#�G���/� ��`& �(�U�ʔ�&T��q�.�����o0�^���_�l$��K��tHS~��zt�S��p�]".��	[�/��g���b~-cu(��=I[�>�.�v6Ny�f9�3(���`,�cR�ke/���������N��*���<D��>oL�X����*u�N~�	�cJ�� d��||���
#��iX`�sp��rT�$/��&��v��V�	�%�&Ը�~ɄD�%O8�_?�z�S!i��y�w���uLI�9N4.7E7mB�B�;_�t�9�V�eq��(�y�}C����9a���)\��l�#{�����+?�7�+��V��Y���-���y������x0�q|�vO�F˨j����;�(Ʋs�Z����w1��`1��[�b���Ѻ����LO�r|�����h3�P�ᜈ8�i�%��/qk���R�V5�I�b�+�2l:n�q�������NB1f�hY��.��/aϑ�W����tu�xP~m�̊��F�d��n�>\(�[ڮ&��ҷ?R�Vk�j(�2��6w��Wސh�/>a� �S����i<�ߟ|"�α��S����|n#<g��h� �:�:�yh�!f��z�-=C}��WP�����m��T�՟Q�-�;�僝~���>��Z����<Yh��T�]�������6��t����۬g+����o�p�XP>���Ѭ�@;<��zr�m.G=z^�K��ϙP;{����$wg�����6������qx	�.G��.}��=��`c�e�ZL�O��ܓR?�.w�@"��Qh����Q���Í��Yw���gKAt��6��
J�2W4ڤLIy�hÇ>v�N>�B>�7p�u�2p���&<���0N/sX�8�dl�!��A�-`��8%���x���/�!�h��ˌV�f�y5��c���``ǀ�C�c=��_^.~(���6�>	PB�"\�X�5�;������p�e��r9t�_^���t7n�e�B�#��Q��3 �q��$��t�����I�ʻ؁�.q��~��3rJkj���;����O
BkVA{ד?3�~T�m[�db�6��U�'�����a]-d8�Âkf�G�d+$V�Q�����Af@�D4��j�(cH��,�}e��?00y.�˳�'SÏdU�P�V	$����� Yx� /n���|[|�a��ɣ�h���%i1����#9�����ɇcwe���)��wݜ�)�{4�&�h�	�fd)m�K���7�p}���ۘE�5�Dk�ӝ{gF�6�{k�S$�����s��_��\�KI�D�R�<cW%��!"��ѷ����C�kM��׬aǐ�D���#�}5�<RG��_t8�������#�lqPN�|Fw-�Wz�t����8L��{�����i��w2����kTT�#�S;/�/`�J�؅?��W j�]:��LZ}[����X���f(l�,y&JK��N%ߺD�V^O�5��^o�6o�+�<y
�0��ַ�ɫ�J��:�x�*+҅�7י�]�~۽��{��ʎ���M��sZNWt��u_�oc¼�R��;���M��e����51]/���B���xX>�oЌ��]\�����I�.��Z��p���Ɍ+~sB���[�ZS�`��g��'�23�.�W�	�L�:��8���x�UA�-���
��
�V�����T��\��O�g���^��U��.�e���xT3{Ԑ��c�M֜�}�ip�W1Z{4�G{���2�����-���,u��A#�2�3}f�ۇ�n=���q�i���b#��B*��Oݱ�4)��vKjY���j��qħl��`*'�W�)>��w��=H��VO���}&d���v,�Y�j��+g�T�/��=!`���m"�g^%���j*g�Gw�1�o(]����R�<)|��J�Ξ�涣k7�����(mrK~�Uq�Q?uМ����
��*��E��9E��!���'���gv�1cP���6����g��v�u���~�l��DH���e�[� ��pٟ�'&&\A���	��7��}yyU�!Ls�&?�0#=$$wh��S_����p� q�� ���oU�OG��}�eh|^ac���%h������]�Ǧg��w�B.��yА�3���,����C���26@1i X���]�:�����s«� L��!	i�W@+��l����aj�q��\OX����mr�q5F��@�ە� #u�$&�/q�Є3:�A���a�I��`%��"�����uLk*�qSSJL/��x�xͧ�F�i_2@�]9��^h����p����#��E��F��&��Mw�!�X�;(�֨&�x�Vq�+R(�U������Kd@d�=�ŉ�����MC���q�e�n��z��� C�x��ލU�2QCfx�e�Ɨ׵9��,֌u�9-�:k,�i�rps}\n1$R�S̈}D7D��@����kq%�y�㬞��Ծm�X�pH�;O��L���p�T L/hcV#	�ߧ�*m�̾H|��@�N�ʧ�����hp�9$�KL��%���F�*��L0X`� |o+_��16GMOxV<"%� �t [2�x���_��!:'''��Y�
P�mg]aT�qX(H)�����^������{Q�o��2)x's��u/:<0J�IK%>Bs�L�%2��7�!��6	~���?��r�,+!�x��ZN�W1���L�B�kx����nX�U|
~�]�P�Љ��F(O�k�)�`�؛��j�l�K~����D��A�x3f�]���R6v�r�VC��vm1�u��-��^ �;���,���\l``��`�iwq[Z���R�$	I(�@˃CCC? $�9����+ݠ;�Kh�I�V��!1I�e��x,�}y�Z]��Ɛږ;駆�p��w� 	Mq���aE����w��ҨG�Xb̤djp>
�~ʨ�N���~Z1�6e��f�ޱ4�y����{���*�LC7Yb,�5�#Xo&H���븰D���h'`q�%8����2��l+9##�Y�]�6���u�@��/�En�A:T��Ʒ�p!Ȣ��ܢl�j!���ե\���8b��ea���E�m��R��$\o����_���� ��7�YI�J�N��$�W��M4-�iSp=�˅��n
�	rKQ��y�z��j�����f�/��r@�f��.�'HrF\){2��uŢd؁��sؽĒ��NFwf�|e���z�xЌ'�K$��B�����>����WJ�~h��i�c-
���I�5gެU(N��������
W����g�K��B_U�]���F��ש>��4�g��b���]¬�Ĭ��h���~�DI �� ��p�S�Hh�;|y���禯�JR�9$4i�\�!�\�x?>�hnNa�{|�Xo������r���O��B(>UK�qH�&���a���52>z�gr�I2H����k	�ח��+x d:����	������
�,K:_�r��L�-x2�Zz��O)�r�AX�&�;���X/�]@��!���Ր�*
4�X��������L�P:�pr ��䰦|qf���ъ�\.���gC�i`\ L>���K��p��:�/�D	�Ĝj�)���ˑ����������ɧT�׫����f6&c��+W�nC�@F�<ÏE@�-�vV�wNӑ.���_�Vg��l���X�KĊ�"��@�g��'���x���^�&	k�c�U�Zcϐ1��N8�׃���	�Y5/&s܉���Gm�/�ˁO`,"���w7��Trm�7�1��m^%FO8��7�1+U}i���Py���T��ɜ&C'K����>)�3��毟�P�a�}�U��R��H��;�?��C�0��x0�hO>&AY�q[�--E������ޥSm����f}���?~� �dn���K�9�������P��/Ep!��2�� ��PQc�Ayn�����L C�{�ӫ�n�:�O� )ܳ*l��p��R({7�	��Ҭ�������ȅ���?1t����8 [�5����w b���N���e����ٝU��
����~oeL�k 䌒h�i�]G';�����{��7l#�xJ�B�e��f-���kA���pN+�J'f��4���C�! #��"�D���ma�:Uy�Թ��zb����p�A0v�v�3ڂLVh�PWBx���MKq�\�[����=���s����^�皤e"�?��j��TꜪ�|��+��G������_CZ�Wgg�J����1 ]C&��O��G���bj��p� �9�/��OB��AHƽ���L;�=��z��˗/��ÕjZG�wɱ����h�qx;�K���A0�ղ8��L�[�fOO�Nfs_ܻ�D
���-���X�_=���@ZX�-�[�%��؜� Cc�Ȉ�l��t"���r�v�K��q���duN�Efյ�m����V��JjQ(J���H����!����O2���zUzD3��XQ&*�"�lR��UK_�/(���� ��X�aط�YG�K[ׅw��O�,�"� �E���䊧DI��bE�3�����7�7Y!� g�oS�z�"���#u�����J����f"����`3�zK[�&I�Lk�J2BQ�ۀ�Y�����,��s?��o;28������aH�4�}����Kh�jE�Jc+cZx=FH�����Bb/wat�zӏ����d��L���8Ѕ�z}�X���͇�.(�� W�y��q��`T�lY�����
�IԒo�3�a�0�����{��S��V�_Ǳ9�/��,B��v�6�2��x�MBy׷=�����	؄2�	!Sw͜1N����܄_,ÎU?>��4��`dsAE.�L�N���O�)��O�%=��=k�9%_r�哂�e��;��,x����,)sss�Uf�d����jU�UF��`@�����]�f����6���5�y#� �����+)�Rnܩ�����\���*�mS98���8�������dA��󤍡[��ҽ�
H�Lww�)�C@q8��(��d!�r�f��]{,�PN�M�q�_%���>}�̘�'M�>�!��D`c��q�i{��vG f~��
���	!|:ʄ�){�\ f��h&i��D�$"�N&�k(�*5�eI�A��m%�&Z�oƷ��/Q������3Y��kZ`��a�hY�����ǩ�%���m`�u��G�:;�x��hl]���f��ꂡ�����B�\v��|���9�m
 s���aLC�!l$n�Z�k ����j�2��b��3��	�ߕ{\��T�WA����Q�g>�.�=�Oa�\@;�j!�HS�h	V����'��%=�xn���4�,ib�@ �M^�[�}�˽�J��8�]��������	 ڀR����_��$+����U�ɤ^O��
O�Xx"=�ֈ�%r�[�M��j��ZB���r� R���61�:��a7:���D� oS"�˦G�}����%��'�؆�fUgF�m�y
��K~���X���+B�2�IW�f=�
���F<��H�6~��E[�|&���p�+�9��h�]p�?�C����[+.�	C�@�nA��Kr*VIǫ�$F���vK%>�ןΩ�1��?�kM������9I�t�������/� �i0�cF���[g��� �_�x����Hֳ7`Q]��YH?=�t�C՜��}UA��Ц�N�Hw������I��9��N.������X��u�Ƃ5n��`��&-��<����+��\�G��
E$�c.�e��㋚������w2���QQF�;_�:��b=ۉp$nB�n���bI�$�-޿K�����L|�N�'(֚���v�������V?�5��(Uժv���b�Ӯރ�ܡ'��B�{*i�jR4���+$r+�?@���N��������\���A�r�;=� ���hZ�-���&"Vz�����腓&���(�M�n`�\.@@d�2yYԣ��c�־��
e3���+R /~sl:��VȲ�}�{����rv�D�ba?��9����c�I���!�^�m������Y�}�~����	�4�Y�(�#�Q�1��!gvp���閌���'�m�RsMJ<I��}v�HJ4x�!�c�:.�?/��tLమ���?�_8��c�n��:�!����lNg��y�Q!Ό�#�����%��4�ϯ �V6-�~��g��FJī�j!bxօca���P�`���l��>{PNO�3��DBMc '_�d� ��8��?b҃������&���ύ뙋1���?����GD"��C�J�!jhy���b��{h�o�Yb2H�U%������Q�y�Q��p�+2�hl��Y�9������ݨV�0�pF�ǝ<� ��#�m)�0{䝔��v��4![A\���z�6���	��/��N5"�zt*\HM�p-o9-��\������ ΅	_=W�40���RɍB�7w�A`�t���JQZ��҇X؋S`��0��ӆE��/ɐ~���o� �eF�r�ɿ��k�ZhX[�l?N�b�	5Z��v��?@��*9�h���(�x��(81u_ !+º���J�h�����7Y� ���H�Q��J�$��^�=*�����\�W�  �몞�cy"� oP���W.�Pq��i���P09 ��v��$|�ގNJ��HҨ{T��~��"�f�I��Z��p��ć�M��x3s�H�����?5$�0ݟ�1�_�x�3���lh\��4�
었=j���0*'s��j��v���C���a_h�t1Tq�wzp/�t�U����X_6�2��r���o�C� ��>]���9�Ӓ��R"��Ȅ��E����HJ^��v=R��@��<�m�Қʻ��v!%��g�����%[/|��s���>��Jv�dh�ε���ĵ��&��'�?Qhz8*�|^�Gk �XHE0��E�BQ���?j��^%�D��|��}�_����Wټ'�W��5�y�䓫����o�-���p���_?�<� r�E���)�`q`u���1�8�PM�lG��H�C0��J��
@#�^v(P��"�����t��.C�b0\٥���{�^x�E樭�d~%$�*ʆ�1�o8�����	�待�FB������(��Lֳ���̅��eq���3��=*~
{��i��
 �I.74J¢�Ķ�}��*]�d�	9Iǂ1s"]�,��ג�Ǽ�J�2P�4�:h���o-4�־ѽ��i���1Z&d�7�;���.�=nZ�g7q��]U��F%!K��na
�ؖ���4p5Q��bΣ��e��χǱJZ"�s�.�"M�C����P%�k�xy������i�:򐢒�&�y�`��m,0��mM���o�-��b�5zZ�/H�ns��A�%������P�*c|?#N�3��G1=��Ȑpi{�l�c#���dRȝm���<���$��cmwUN{�CA{���U�X�wcB��|�A14�˭����Fp*$d�1�r3^��<�������gDu��WH,�}��]��}u>.�Y,��������s��fa�b������@�s\�>��ԩ�[�~_�A�q������4���jf�H3��[��"gY�K�ƟH�u��K��%�"�Kv@`���"뉜��R-2��yD&wSUd�Wd�,}���j�W�j6�N͎���G��8���5�x";�� }#<Z|8g6�L��{��ލId�^ͻO
hi8i߽���_�a�Ɯ�psf:�[�+2�4v�29�����m�։�V8a4�{&�W_k�7שN=]e0Z��Z�F���vR���O���y�����JB��$le�5��x%�P�����z�\��G���U"r��;�{@�����((�@\�Ap�v�&@
W�o������^�Z-����1i 5�����)CՅ�fm�|��%qr�c�]�Ľ����YtZ���<Т����� �@�:�T@����U�D��L�u��6ߞ&o�Љӏ��`>��HP�'�R�L�4����cp�tt���-��tP�1�8��ri�V�ҥt�'�q2�#�?0�
���B�I�= !='�]����{�r|<Y��_�蹦l�D~o+Aɖ�dZ�E\.X���'�U�o][`����w�*8/��>`�a�w��vj�ec:K;nO����O�^��%��	�g��΀���d��:�0����2��Pk�]��X/{4x�צ�]��й�\��W?�� �W�bvp�_zI�";kv��6�C� �B�������p(g�F��h���/��J�U1�����J��h�- ��[Λ�P(��Z����s�r���;r-2�-���	����t6ΞE�%Qyڻ�:**�G����	�����dm�e�ÿE�C���|>`��s�[��/3�輾PGEw���[��q�uutpO�N?H�]���E�S����ɖt��ыc�ٔm��)ؖUc3��OI������y<U��~��B�R�LE�S�DQ)���Ǎ�*$��
ɔ�c	J汤c<�y�=k�sNw������{�>����Y{���������{��诎,�jLU��	>O��͝D�B�}�}L�У��H�O��K�z�Xl�~���K�����؆O�M�R����.h"�~��+�t�H 
��#��?\1gH�B��
�v�	��8�V����T����.+D��W�v�H���]S������q�����A�e�4����؂�OH@�����ja��\Օ���>��D�f�s��e��9
��H�fS���x�I�(K�c��S)#��(c��3<�RP�t;d�ݦw�~Zm��p��P�L�V���c�!v�>������k2؅�y@!c�ߟ�ֻM*J�!���k>]?xG�$K����A�cZ+�A7��`��@bO4U ��|�^\�h�ƕ�I���un���q>G��##죜e.��~���q�uGvb�_�J����������X�腤#q�R�<==��� �	|��\8?�(Sr�Uׅ���C�g��{Ze���&�Un��>��eР#p݇1F��Z1�"i��)�p+ܚ�6�vni�kE}#P�X�BS'\ʶ
<��gP���Y�m���P�\�l-)7��{nB��j0	�����W7�d��\P�.""R�� C��{|��nT�M���l�ٽڢ���I'�Y	
���i�h^�ؑ酥Jߋ
y5FZ��Np_���8u���t�5�&"��*#�\jv0l�ĮU�kw[3�H���s=��Tm<a=�QQAS���ǋ��Qh��|X�߬���������U�ݕy��f�xC	>��؇hL��j9֐�n>� V&��!9����5׿�){g�&�dV29���X�^�����V[,�{��n)����X�)�U�5��t�ITo����m�[���s`J�&��F�z$�s��mj��::�v���Ô��nh{�f���[3�J�\�в�Ǐw�r������j�`�)�䉈��Hu�oE��Y&`�V��e+'Q�� ��a��xܟ�g]ݶ�\D=��y,/�-h������|���h��r��e?� YC�[�\�C�vb%���b�ׁR��N�w�$Wk��
�t��_�P:�u��� Uc�0�ᶰ�l�O��v�沾�5�P8�\{h@�Vq�F-�cbb"�, �k��
�ek�/��/Wc�tU����������kzǾK�LSZS���J�%�Ã�b��F��;���x�F�����Q����Bh���zbh�!�]������t�EH��E+	�[+����	�`C�t��D.g��Z.F�Q�8Z[��o�n�2�.�{/�A|��^�#ga�I��

�(�9���%�0V|{��T��z�D��_O�F�pd�ۑ$�ؠc�K��}�����@bJ�����\|e��]�����A�^�뼗"��1��������u�7�˿)�3�S��*�6jD��r�W�<�
���;c���=%Z�<���"qX_P$Ol(�M�>k�-�#ia�0��l���0F҄��%Rm�B��*Bw�f4�J&�i^�;�R��i�7+IU�a3<ʝ��"d�D�3h��&��±����M��s���ۀ)ڤ�9^��'�������e�=��76|b���*Ci����W�AO��=�߳��e�3,�vx;>�3���鼑g��G�?�}>|6@�1Ä0, ��J	n�M<���h��gAm��ryA�B\�0,!^�+��l��/!Hێ��<Ӭt�Xs�#�U�]�ᙅ
@u�T*z�a��8ĺ���Jx������f_����%Q�l_��M�,,u��f�bg�3���Sw,Pu��J2���Ų��?�b����M�a����d�\R6�+Gy��J��ZAsY`I�H�q�cn:�I<��|��w+�E]���<�~�8{?f�؇|^(��o�i�Q�����־[\��h���wg�ʥHi����7���9ԁ�[� ��Mc!1�{j9��!_��9;���,ļ�A�����(
�t/մ���ev!��b����ٝ�(:�iJ��o2��e ��c!z�l�]���V����R�æfH���IG��Dm[wY�	�H����EO놓�f(���l�-��v��,Um������C�4$}ꤌ�b�>���Ƃ��XO9��%���@�W!V���eQ��u^�4@g��1�@�a=C��``g¥l�MX�U�E��+k��:B>=
�����g�q�I�w���&$���X0�G$?�q�b�ޅ��i�-��28j�� ���$����| �́��5�Eb�(�:�}ؾ%����
Q65� �chF.�ŋ�oC���	r(��\��<ע��C���v<mE �j)�?�&��8H���	J�[�X��=i���P�]��w�0d�:��Lĕ�=������7�I?����
�Ny�s5ٮ*��AW���hP���2Ԓ�M#��T]�5WW
�^U���e
cn��F(�C��)�s�	h\ߧ�;�<�$;C�P�I�oͦ; �I�^>�|�᱇c���̡O;�
��Z/�h�����d]0q���G�G��L�)u�=YP ������[��{�g���z��X�]��$y�m��P�߭h���Y�U�t#z���f���e��;��\7�j��5�*�_M�(��[�$�T)g8k���*.��b6�"��^��:,�ZN���F�� $>���@q��5RK��gKw�@RC�/^����o2�������G��}M �J�� )��a�)��M�����ITfmD��I=������2����J���˳��}�ɶ��|�A]�t"U1��z���0��@���T�S����z=_{R�鱚�4�����;#�
�9A>�ѣ $���c��l!�O{����%0���-r�Pi��I���b� }���3q��!`��h��ᑑ�i��^�:�0�Զa��L��|��܄a�o��+�{0�;�E��b��$g<�w�S��e��L�L���:hՄ����M�ô)7vz��c��$LmZ)�2�F��|��,��SFn{9���(�A�{A�S<�.M;	�G0Y?;!�A�F��RKɁ}�ss92G	D3GVEA6�^���XIr��S,ĎH�����_�J�Q��ps`��u7��V
��u?�A��<�$���>���:�6�r��|II���b'g~'�0P�J�����p�����A�ډ	
��5U�E��gwm����Hܲ���mj�b�QzpF))�X��D��,$�xQ�>�/%u8O,�M��	}X"�}�����!]IHTE��I;��u_C�ڈ�{T �Vo�lC�X"[��Hq�K�jp����I�&d3C��I����z����1�޴�/5u�.�V�篠d5���4����{*��f`\-��̩}e��P,�Ӭ��jT99B�J���HC_sqNO�P�Px�=\T�����#�s�Ά	Yp+��S�L��J0V��H���q�,�����:@rn߼����+�[M}5Y�f�5�D3,���2��f/��Ր �>r�t ������BII��wP�� �Ky��E!�gx9(/�2�|�� �ěE�x�(�PN%�QN�:Μ�W!�,9�62C��,V�Qd
,�����_p�r�Iʯ�Z��#���|Oa��Ơcz��Ux[q�~9D�E�����*nSmc�c�ވbe�M�RJ�c`� ܨ@-�6��!a��M4�܄"�pC)`�� +\�#�{"��J��`��C1줪� %Y�w5>�"�s`��|F�Y=�`U�J�v��s��D�^�x�{�/��IQQ���s�9�"ŭ̥hBkV	�@�fv�w ���-b���WQo����:8Iυ^C�9i.��?!X������ÕJ�V>��HsqW9T(��:����.��%�0\��>�Ts>���6T3�hZEp�Wx:�x���cG$}��b<>:��GK��.񣾞�O�8��V�N��HJ�_�^����<)buސ�!p��Iw�3(����Y�B� JI�C�9M@Up鉭%[���e����Ao!I%��ډ7բ,"�>R;�I(�r��W�������s��)hIBVb�ɢl��#74����}�Y���D��jj���5��WcU�U��TT��9�p�MX����.Fj�P�}��l�����e����'PAck�H5F���8���舢U��O��Z���Pt7FM����q�M�R��}t/��6ˢ��M�b3���p)�xs�����t'Z�g��@l�(�hM߶���znL�b�麅�S��������#�2e�0i�L�&<*RW�����NM�UXq]��R<��ϔ���&�;>M�)h�K��c���Y+�8��Cl���.Q�`�xG��\F
f�4�]%7����L����˛��چ��N���UG kB�*������2���Xj�v|-���ީ�w>K�@��H|�2��1́o��Q����m?�s��nBxz�|��|��b理5k�a��[pSs�����#8�A�'7�t6�=Z/(����M`T����z�ގ$9B2$�Am����)o�ȱ%�a�ނ���M�%���1jU�.s�@��F�&�� ����1��|Jb=�0����A)Z8�
�k֨
�P�ƶ�"9Z�f��T��\�T ��0�M�be.V�R�.
��rz�%8A���C�WX�Z�WJ�P$Bqkv�	��5d��|BoB(�2��N!�HL̡*�����!{��H~�G�C?��pގ�,9��	_��V^M���n�8!���@��3��j N�t�`�'P>�TY�Pi�޲>�̈́�m�0�d��"yxA�44�YF�}7��wʺ��. ���~C6`��<
@b�.Y�W\�̡NFD��j��x��g+�zPF���	Q��ԙ�0�f�HS{%�\�E(VE(c�R�s�~(�\r�����+��O���9���T����Ji0X3����$i���@�"����GsHWX[�B5Zoۆ]7�\�$�Yyz�{to�������*	��x����"u�����C���aX�V���PMa��Bf�cᕷۉb(&|"��|� ;�cMD�ɵ��7���#5:ٚK!��1֨m�1�y�C�Л@E�/ �;���#M4��3�S�&dG�HM����qZ��{4��܃z||�w��Թ��z�I�Gb���o8�(��2q<L�s��c�����̫ E���"՘��^
�P	��赇ˇ������/��G��#v��ǃ/�o������xmZL�P�#��ky���3�j* ����ԃ��Tc���E��k�W|e}]k�E�e�4#�M�B*��H��O�Me E!��ԸXsg_l_� 2F�n"	��Jȫ�65>�ʀ�h����o�%��4�N~��ޢ:�n�h�P�����s���w ��WJQ�Ձ$��JGٌ���<��� �7�a͜������A��X=S�n� ��x��s��c��[�sC�ч���>����V%Si>(xΎ'^��*��(�ؾ�qtޤ���:���y��7A6�Gq�N�"�ɯYnή_�)�FC�6>k��U��+
��Zl|����U����ʐ#6��L ��Ύ��cZ�K���"i��ƍ���!��gkW�����M 1�^��n��m��z��V��56�mH��l�Y�w��6=�����Xߛ������-��y N�q�w:������X�P �v��#4Ҿϻ�k|^��S$��2��7(s�F�8?��d����A7P]T\E�-���g����2Hӆ:��5-��CS�B��W챬����צI=�u�s5!�����{�2�`��̲l��+�A4}�?+A�k��)d~�����v@��c�S�G����MWs���d���~_��eÁ����F0��kf�vr[�Ү'_��}u��������{ʴӐ����Ⱦ��k��?�X���
Y�KF�<2�Z#��u+����ւ;�m�����u����@��HSEČ@�.�و�\�?�3��h����н��U�?*e*�"�:/��,O�^M ��r�&�Q_�'n\{�O_b���bv7���#J5FHa����Ѱ�����Ԁ�&o�|�*���n=�܎�3�D	�G�������~�ߏ��~$�Tu(���8D�-�OmZ}ZcO��⺇t��8��"�OQM󋟌MU����h���X����]=zϘ���4~�?�u��ٛ{�����M<��hQ��%�U�Q��pt�ӾضsDj�#Ƶ�_�!��gb���+�*��wq�l�����]7���^���������]��K�?si�i��˧�������ePr�ˎ�X�KHNNVB�Y��W��P�h�0k����Ǩ�*�&JYu�F:�OՏN^W�T�bR���i�_F���C����U"�Ý.��o�R��o��,F��<59�>88�pN(��1���(��7�y�{ү����b/����ܻwϽ��C�;C<뺁��M9αƞ<y����´L����j�&����&���G]\\�ǀF[h�������0p�jp�t���je�Y���9���%E!jq����h?�H�Ύv�V�_<������纵k׺gx�,{��Nu�J�;R&����>n%-/�E��¯���P��w��o˼]u{������Jzzz7��f�n߾=�ۗ���o�98$M��uݾyS�z�ȯ�+�ʦ�~Qu�P��PTM�ի��z۬���c����n�9M�V~aȻ�[qʯ!����r�)����J��1�@�^��]����7�Z.�u������v����٠
���և�e�D���	=�{��y(+j&���ye�|���c�jWW��ٲ�h��jv�o�d�R�D�Z��!w,X`n3=I��膍����e^)���K����hR>���͝�����[�edh�)�`^�;�{���ܖei(c?�5�P�A���i����j9�p��h��4�7��$��������]>h��)��7���r��`����L*Ev���7b��e �ˮ??�u���c��0=��<J��kK�y���;Ff'��8���;��J>���/�n��u�K:�\%�T���V~�E��Ƥغ��n���aq�Q�量+1�"#���f�>�����
��m���s��Ϛ2�p���b��c��)������C���
��s�g���Mz�f�����v��H��)��8+�����#��Z����22.5���z"!�eee��UW��kփK3]�t_�"##=$�gc븽G�߇zzz�<S����S �'Qko�i�� ��o>+&	Z��v,{α��SVV��E7�<;;��B`��Q]f��t�;��������xw����2ه4�!�+�
�(���T�hh�<������	---3#]
[s�k����k��������Mj��#�@��`��촴���X1hD`�!�[�ܗ�Ә�EˆGM�K��ι��IۡX�*ܫ��iCGG��f�&�fv����˗/7�/��Ɏ�����>�k��]=Š`��p�ެ�'���'��+o2�[G�}�����L����{{�<��^���Xl�e��2ao��������G��E��JQHH���������p�J��ğ��K���t� P���'jZ�M<��|��m�7���&�QU��: ���Xؘni�u�Б#S�?~�������ӨE����8T4k�u�֒X��Pd�V@�d�-��hg]��Rs�Qy����G^���`����@���הEB\���e����=O8th"�"P�<�͡U��\�����S~���ﲲ,�Y�,uy�**ZQbbƈi��ĎvHF�����69�s��8�U�h�Y<".&6� � ӋLP��k���k7y����RXX(��³h�Ql4�mB��]�����d��ڙ�[2�۫��D;�<V�������9W�v�����.8:� �t%��WɹL�r`u �.!�p4x�l.��Fw�������J�9���W=:���/5�Bwz����`:ˑ�<G1;&?#��8 ��mxg8�~t+����L����Ǟ/����mg>s�l��x�<�Uo�os�C����C�l���)0��Ç�W���gQB�JQ=�G �M+,��6ض޻#F/����e��\歙 �u�� dT�#��7lX���#���oL�S=v��!�0��K�Di������|���煃U\�xLO6�ʰ�v�*��T,0J�n���=�W���i�egg'g�1S�<��K<\\���AXZU|��GEna6_�}ripp�iuu��>����ѡIo�=��������障�Q��#�%iu%7%ed�t\�5�SB��ϫ��.���c��Q�c���'�w���FejldddГ�\��B�YqF��c�������]_�%�<�O��HH�m���|���I�\���KGr��]`�j����7o�p1y�D�MG�e`�"GKmdf^���s������Xڱ�no�!V���GTw�h���r!�e=q.(��s�(���E�'&�w~����xl�8j��ó�WSSӆ!|�M�wt�~�����LLL(�����~Ѣ��N-HU3h���pp?�/"��T�;#J����@.�<ݯ�Fq	4�RRo��y+]u�c��|=�Eb���,���ڦ/-/-X�(<���T���c^����vL�9����� .�@�1arp� �1vƼn�e|�귺O��x�j�d頗ͽ��k��8�z��)�oV���ǼsNZZ�ѷ��~�ɣae��+�?�o���o`�����M �	d�U���3[[�Z����3���(e��ny{�ܞc;B$�XV1?0MN���PoJ���=:�Ou��)jX�x���xRr���S��mFV�6Rnab�7F�{�d$J�i���T�xo�zmr�B��Hs����1.�rVg���1H�ēv����,��C��=z��FGG�@x����\U!�y�0��q��Mr��	8��Z����^�EǼs��Pe�)��O(XH0�����#e�k"dt���_"�y��x `	/v�b��))�SM�tMm-���ٱh����u@� �C�Qy�� �ۏ�3�����8���71,y�����yh�ܗ��׆��xO???s�^��Ml}��h�d�]�H����l{2���^d�R�:�3��Hn驩V��Ư�4����"����-� �ج�kןx����Ex���o%>#��=�3\fȱ k��1�R{<��`��<�WYY�\���>�ݻI�V�.�-VKRT=�P+wssS�����x����Gx����X"�|����b�$��$���v}�������	Z����{0V�s��e��U	d��|�1��/J�a:&{o,��@�E$d��4!g��y��V ���y����۱�222�A�T���Ŭ8@A q���@�34��w=�I.�W��n9��q�<t=Tm�"�Κ"!z��S�����':�tXǭ!�޽���#+�KeJ��'�G�<G�XqA0/�́�Y�<G��H2����r갧�'��Ĥ����z��#����@<���� ����N�/C)f���" ��Jq�g��メ(�d������Vb�' �(��Ub���2�J���ۻwo!T��<��
��[���y1Ӳ�}xB�L�&�xoN	�|'P�+G�Ubq��C[����Qtӽ|�;*/^�ݩ� ����qȎ���}}E�b4&H!R�u
�=�s�'bLٝ��zm�!�� �O���qZj'j��䏲��O�I�T�{��3Ӽe��S衮���]:Ve��[j�
Y����@SR���	�"Y@ˮ�][�Ӿm�� �.�y�իWk%@z�&x�2)i�T�ә�۠�f���g$�tKU`�Ť���ֈjcЪ:}lх�#~J1u�����mPw-� �0�}�Mu
kT�R�Y�\h��E�u�@#V]<:�Yut;x�)��ι����X3��YOp#)����ў�/_&_HlC�V���[��Y��!�r�ܺz�ƍr^�Q�`��.��3����Ʀ���-CiJ1�2vLu�?I$Y�TQ�-?&�� !��@%y�(ݲ�p9�����}���PpΚ	����Z���\&{��kAJ��}ll,뻤�+D-N�<�w�ӓ���1��o�~v�ٓ	Z�[�x���	_�����`6`�4�r�a�<@𛾀�]x�]�.1����յ�T���Qǧ����ʹ�ndԣ�K#|ie���ӧӐ�<��nC�����Y����u
�لKI�@'?�����pI�"Us,��IU�/��0��o��4X��
��n1�D
�#V����0���|g�Ԙgn��Qf^�řr��>��Ǔ�L��ױZ	�f;� G�%D�p�q:�,Hluᐆ��333�����A�VY
�t����h��x^�L4���3����P�Ǩ�K��Zv�_*��NNq���x7s�!@��Y��%��:Յ���"��}��)\�	�h���a�uh�5���i��f��5;a�`ٵ�9�1�N��״��H$?���9矟B����^x@U݂���wɚ+������ӧI���:9�J(���
'W�Å�:����Әx�A�h��}��i�1�������~�����_�Y�.!v�Uf�}�V������d���� dO7��:͎~C4��h(_A�ӧl�;>|���j��!Ë�*���Y��7o��p6C��{&%@h��@��z]�K`CI��?��$%%m���6?5�lٙ?g��E��p�a��I�G����)ÞK�}���[./''GƎaSH,�p�O���8��Y��!��s�,J�{%�PQ�Wh2B��@��l �IOCB���c���dd��jBO��w�t��3�q�^�ڕ�Pub!��d]��А�(��������4�S�>�t,O�{.���̔�u��̂4�fU��Ie啃^L�}�T��8�F�T�� �n]up�.��Q�'X�����Ւa�d�r��|�BO�²1�">���`��Ƣ��q���O�*�^{��`Z@]����?��sƕ���"�����`B�}0KB8��2\S|��Ĕ��m��K �Q�E���J�}���*q�F��nEPT����Cpzh����;�R,ѽt�5��w-�,��i�#o�t��Z#Tn��� Y{k�â�L�|(�)j�xTΝ;���S��ꬥ�X��������&
�<+K�Ss!Ե�������a��pLB}�^Ksډ�Aĸs��*��U�4�?���5��m�ʴ;]���󈄄�^�����b�XO��7�=���>x{�	�F���[z'�jA�������9�>b�o�=��n�b�U
©�Gr�C�t3��pJ��p�( ������J
qm�/��Tz�Pqkkk$���&)�;�~��Fvd�����A-h��\^*�>�7�yeif��ƍ^'|��˘_�����H\\\ d��1.%$5�ne�n����3Š`@�?����c Z��.���2R �������0__�q�K{{{��O��EF"�=����{&��3�$-!T�;I���&�?|�(X������^��t|yߠx�e�Ͱ礝�� #a��djj*if��C�����S�ez�E�ҥ� �c9�d?���b<�:xZ�;?>��M�A{ɪE&��jj;:���/�̸4���ÞIzYjQ2�d����;��hW��L eY� �;_�����]K��!�wbN��ؘʈٳ`Y� �P�����*���;??��2��������}��˘�z@��V���/�t*.5����aO9 i.���5�رc����ې k/p�r�uk�����v�*#�k��W)�����k i�			=`}��Λ�w�a�߱�A}����*�"��i�u�3,*ߗZ����J��y��`���^# ��)�9hpS�J��pZ��|sf��\\�ӝ.�H)}�������EX}��t�UUUh��69�F����}��90n?s���da����#h�Q܎髒|���lO@���1�wGa���˗/� ��%pR2]}��!C��[��8Հ�l��"U����ðv�{]}��(t�h�	���]�^�����Ӄ
��4��R��r��nk�,�9@Ƞu�!��N|~Z�]�u����R<���ۄ�'���1V>!���}�L���w�����K�7�-�ɍ*��P��T�v�^���R���r҈����{�%4��E3̞���(��MɗexO���qr�oh\�ʓe�������`���i������u�[�QSu��>r�Mo��*�>bڒ�8pl(�v������C&P�"�٣$H��c���L Ä�{&A�����	��*�����R
��&���B@�h���]���Py�;��Q��Xc���%>,�]>|�U�x���_��"������
�� �B��~���&U{m����s���}||VD'C�^ e�G~~��&�u�%e[�Q����J�����Zu7���~������m!��z��#E+��B�6(���C�IR��V��[WAȡ�� k� H��22n�e�5��/_4��V�_bEkjj"��$Yi#$�n]��&)A4j�Zʲ�ZV����y�@ᮡ��/8A}����I�1�}� ���Zl%�X����FX�@�Nk�x����B�^�vP�8���M��F���e�.��)?�=gBK!y�K�W�ሶة#;s�l�>6��OȨol̔�z3	���4p�4�V�"&]$�}0{�~B�ID�'<2R�R�V�����FzK���f�C����p0��|E W'�U�C��#G�H�&�P�Y�_�����O������)��>F���?�#0�[� K�ד{�>ntt���Z]��]�F<8]��(z[ \$jaa1��"�% TP3���kkGB�ސN���/��)�]�
ɦ������@��*�:��6Te=�%�(��a�%�=V԰�U�n�F�.)���7lX����׾���GKX�.&hIS���k�*�������	��a��ӷ2?Nz�)�vC322D���1�����n��ǃ(ϣ}�������".����� ����H?��,����*g��G6�����/���p�����-3jt�h�c�1h���X���K���I?N���a/�*�ہ��3��sn���[ɾ"s?�G�鑳mvyc��`ڞ��Q�=�Wֽ���g�Pr�|:���kF�Ɋ�*�n��*���Bz����{�y�`�.--E�����K�H;�(~��K�+I�j�1�疙v i��*�>��e �c?~��[ �^�푔:t(���f���Y0Hc#/�7�>�+nz���QϞ͞p��VR����V�Q�7���x����q3����q��g���"!����
��JrpK]�XM�%PtK7Q�yí�L+���󰰔i0�;�S�IY���@�qǰ/ә�`����0��6��GY�LȦ�c9��
�a���~ժ�����;P�)�z�
+�)��P�~04�SmmV7�Y�]`��`bb2��[��U�r��iZB���k�����ڳ�@��=v�d��ͭK5V�q�|��Ғ!�V��
\]�2$���..�N է���a�&w�ܩ��@*�1�S�"�gH�� q?�k�`�m�N~C�͵Cy��3��Y�_A6��Oqh�<ZKHۛL�3<�x�����$����\&�9ϟ?�+((����I��T�cǎ��������<R��>QѦ���, -�U������\�3>�9�;�i�eC�v�8=��tD���@���NW�!T�ǕC�	��~P(�(�����������N�: '��6q��y��e ;!C���Ψkh��IK��c�� j����ɩ=Op��c�r%���ƾ��G�W�)�
�A��o߾ՂM?쀄��Uei�Kp������#G���H5�������Beb�!�Z^Z�C��}),,��GS���xlI5q`���.�N��N��?�8� ��`��H!;L�*Ctw�I5�%�(���k�	sgA��V)���6ʳldm��`.1 u��x����Ւ�{�2^M���^��3���LM�nD	 ���+�:5vw/��l�*���s��M�k`�<)�M)Q�6.0�}�6?�b�t�9����82�un|�Z�.'&�)�/�������p�y�LzL��ń��,h\��l�'�ړ�ݷ������ݻ��J��QQ㧰b����Y���4T��kiӭfQ���A_K7�-�vY�
o 0�b(oo�yOOO�sہ<��/�>��"#%u���^;BX9H�y��������Gt�N!�F�M��B��&G�,��`/\�_q�v���/\�p���< ||E~��1::�~L�`f�抃�ە|9o�����n�&P�� �B�WU��%�7"(�����O��6�?}�����v��H���J��Rrr�""##y}�D���~>,�d���}ڔ���q
R=]�O�`\˾��50ۍm��}P�D�W\]�Q��K/5X���V\_���
v��ʒ����j �j��
�x�!,�j Ԥa�Ȁ��uu��h�蕦ࠃx���-�S��5���L����[�#G���!=���+¯��� �
�bS%�i�;	Tj�ּQ���J#�0�q��pGggghB%
��ADMS��N��@�#��(ds��4���C�8����j|�����t�������MT^B3�q�f���+�p���orjۊ������)�v�q��C#��|��h�7o���1�E����2F����q�~zf�/Z��03E�;��&?�����o�7b�w�V�CM"�o�^�v[uR
���_�"�3�z��kkVF�R_]̱ofO�g��w�+��S ���ˮS�y���\��)O�p=3���r������R���		.�Cs3���n@��dKNɢ��\9�i�i�Q&��{�Ϧ�U_D'��AiB�2V��RٓgϞ=���A:�>���Xȃr8�W��:�'|&''��~���R{�y�@9Yx��y1�j����[,>%����~"+A�5+�n' �03;�� �����y���II��s��z{�x\m�rjQ|M���G�._�C�^�}���@P�*H:T�GO8=~��ϑ�LUrs[��,�+��}A�s�m�im7?7���e�^uu�-��-��ݓF��@g	�O���T�����젆� L^�~�G�Z�/�jԅ��GP����_��v�b��!Dۨ[fff�o�^-t����0�\я�C��5�N���n�����B�6�1���;�������Z7� -$�K�L+V��߾�$�8�ف�x9�okF3�A������g{�T^����n�́qJ1��ոl�b���D%�41II'�_�=B�"�;��*D���]Eq�ۖ�D�?�Q�T�_MS��;::V�w�R�0NOa]���h�ny�!a��K}��>6���J�t����%�ʩP�����p��*?�7p��˗/����!;�k�9�#G�a)q��J�}���1h����q��iG�-���E�Ղ6hμ��~��cqqq��]��S�琉
;�����eC������ ��>s�-q�v�=@�O$HF�����B�N'Y��䤝%޴�����d�psZ�KԴ)����s�|$�R�}����:�nq���@��W::�V]���PFVV��i< \e�T���� >���ۨ����S����꾀�----���Ǡ��v G��xRN�,/�,��?gΜ���q�7
�BM8i����-�;���XF���Cg0m ����_��qs���J�!w�\z���s�U$ �e����c��O���]3������I"Eq �f�����Eź�M??�� �}�*1����Pz��9!ʋ:\��,8�r����U�ג����Ԉo~200P���R��6��QI��W��MN��_>�<v��B��ɒ�/��hB�=>f�>�;��QB���ԏOL�K�
�T@�L�`}��H��vmmm&H] eu7�l=��TT��q�v*T���z�_�����$���zB5G��	at��m��1�I��ހW�^�+�M�Ӛ^:�/�ͤ6�a����ܶ�[+�D�+�|����g��ݻw�^�»|����ԓ������m:���C�Ӵ�F�:�R�TfFVʍ��/C}|@\|���!��YXx/������B:�weW���BeaYf=�5mp��f ������o B/�T2�wH:*���q�����}	2��+�䮢��/��$P׃x֖�ar=UFΜc-E�abb�yOb���o����4�X���W���Z*3��V@��[�Z���>F����J��|T�q�h�M�S�k>*E�^mhl�&��rs��K���
�]"���K����Q!|r�[Qz�D���|/�LW���<8�b��Eo�!�SM[��KK������>#E��8���Ń�Ν�iCx`�`v�!��!>�Бwi;�Whc�|�ܷ���޽;���]��(5uuG��'AW����T\O+(X�nll4�{Mރ���}�`����w0�`����zĨ���v��Չұ��]_����������w=ހ����&g�2��*CtF��r�]ži<�G��T��tR�z�t0�[y��Pa��7:TؼQ�t�%:�������uuuU���ZS���Bt��GoUH-;U�#��T12ꩆ����� ���lڈ��43R��+�?yrrr�6 � Ȫ_Y6l�ϥ	��4����ӓi �w�I� �\�{�k��,>=�=�1��m��K	G��
��
p���3�	%E�~;����A���)U��Ă����F��,�1!��
���軪�\�v���)j�oe���q��JG;;�f(�� ��z�>ԋ!P�S|�:`Y�s����IU�*-�3}�E�ݍ���S��i-by����ec�UrЮ�":
�s��Z��3G�� [W(>p8"v>|��ԑ#S�8lü9)�p���>��#��$iǨ�aj�I���5ƴ�5�z^}id�%���1��3P�	�?��W��Cuƻw�C�����T�ct���&.�������ԑ�4������"����:+u;���l^$ltuE�U(��z�����a���P ��;��H�ٯ�OTD�g�<����r�Ǘ�r~�������6%9����h����drS}�h� �;wޛS��ß?�"L�T�׾�O���4��G�؁C�CV����-��x4v���Pg�Ry��A����#�psS�A#SKhj�=ǖ���d�_�-�2u�t���Pe=1wȤ&=0 ix��&6vv�{�X�Ԧ��T�������˗� ̎ ����6���� }%�s:lP�|��O!�`moJ�{����@���J�'=�"^��ᬕ䎼�n"dJKP&7���H�J$y��P|�H�\-aQ��6��<���A��z�O����q�6��Bm��D:j�e�!}X�A�?�άm��ha���q-lhn�m��0���9T�����r�z�gX@���
�}���_`L��[L{گxD��pe��X|�&�q��v��b5��/�UPc�+!9��EJʈ�\ �#22?�,��
��pٝ���z�Z_tg�NH�ikk[p���RA�_\\܊����}��C��Ǡ�07���}"��Tg��Qd�Ӑ��LLHY@�l(P�Z�x�[������yiS^����h���:&!����Y�uӞ���Ԟ-�X�¥�2�ֺ�P��~�_y���kH�T��b�j9��F?	=��=����i;��]��x$+#����͉sA��wX�(�L���c�Ow������g!�(�|V���,��To���ӌʓ���:7n�*.�W���Ϲ̐����6�y�9�s$������H)B�J���-�[�ѮԀ�;ck;�W+7Ӯ�
'$h�ss/��*��� ����t��}~;���	��A�2Ys�̠C�{��(Zg���G'�@KH{=��Ϟ5K��.^�*�ƃ$��6�h*>!�A���<���/4��� �M�͝7�@lhhF �J��R1��6��J���n�,��(�2ɉ�	��̅���q�Sũ�*��!�\n*pE���>syyy���ʩ&�
��o뉘� �W͹���������[��m���~��� O"W�in�Uq�m3-Cð����)���Q8y���V�������������ZI�c�&iq�줤a^fn�I��M#�0����܉6�UIII+�Y�*TB�]�v���a_Z�lx��oL���UP�(F���`H#�� E*�8�k"dj#dfRPw�||jϞ9�x��5x����{�22\����qD+�X���)��/����[��f+�DBq7��+S+���#c��<s�r�(��3{1���ӓ$/�'�22��'��_�A	Jty	��&D�G�4���F
Y�!@̢�w��]{�Ķ6���Lqv��С����;�@��.Q�r3���� DB w���Yj!51��=�*7�ח���rPG�$�߿@^u�`����}^,����A�S��+3�(*���A�Nb�ܱ��f�����k{��(J�{*�*os޽��?�M�J�-y�\<�� v��v��m�\��
��g�����yPCT���-x�8W���J���Z�$�E������֗a��2��'ҟAm��ǩ��$���u=�G:ȸd5�G��"�*K6���-�z�W�NTK�B�i� ��>U����Dn<��J8(��RH�\�92<����(���&��Z����me�󅁔�$:J���{+� e��-"6��Ξ/))����2j�}[�ߒ����?E���J��1j�˞��.J�@�zfӧO�)�jFi-E�����o9�$�j��Q�]����i�/QR�?3�e\A�Vf��j�������`N[�0�z&}�m�����(�Wg|nџ�Z��:��H]�d�ޚ#��S����c�>j�3���/q{e����݈���MI�u�bbii�]��Bs;-z�;\Vz�&�g�L�����������[�Z����0������J���Nc�2�k��#T�ji ���$�]��	Ǒ��u�Th��|�Z@<v�X���磨�e��<������&%��$�M�+�T�8�x�а�Q3AK2��7��4qq��ׯ����n�U�AD���cJ\�5��(?�
���!_����z��U����eō7��]��������=1&�.����倔�8ˌ*P��kkkW��j�R]S#2�΃�k��m��i5*��%ǆ���]٢���M�'��2`�6�9��<��³����`ͯ��Qa*yձ*Yv�ӡ�� �Jm`E��Z�#����WI�����؟���t1q��$M�C�e||<�ҭ!5:��;A�!i��
�YT/��!��S���G&�?��1���l���~-�����<���n�fݨ w����Q����U�<����1�q�z{���}GN�
���U�u�P�0{P����B[=�6ll���(.��Aꈭh�[-�>5�WM&���� ��@=?E]��˲�����̋�_4B�^۔��&Q��TFG��	oI��5Xq��)_W0�	 S�@FB)�?[d��=������ъM��Ѱ�y���G�� e�WT���B9�ҥK�P��&&Q�P�ւyr�qk0S[W���)zzz
�FEy\��uM�5g�b��Ke��� S3�<n�Օ <��U^`}�+=�ߨԣw���q�Ň��Y����`3���j(C������������/�q��ߎs�A��R:�DR�䄢TG��$���ގ�hD�f��4��aG*%�������n��g������|���Ϻ׺ֵ�u?Se� z̲��}M
(^�'�|�
/�έO�����G�0:����Jv�m
���G� �8�C�ƈLU5��TyZ�9��oܿ:�I� ���[[[�n��?�/z��%���Q˂n+3=�����(VU�<,M:��������R����]��ON���%h�"$4]-9=}�/ee������B�F�9y�ض���Q�?���H�Y1�����5�+?��Ĥ��_��]�a��齷��}�(c�m�������ق;���(���T�BU$���� kgi�I*5L�{f��E��弄NA�WVΎ�ܖϨ�9��r��m�!U�T`Z����|�:g����T___���{��%j^5�*�E�f������?�뢱�_�����ϛ:��m��?<��O��o��y�m�c�D�_�w=rR,�HHi�����M���{��3��A-��%�c����G��0i
�u�ɽ�����}�|o;�F�s.�Q�|2T#Q�6"�.q��u/���hH�nlè�Ud	��N�	�s�.������K�-������l�k��~�A�m��[�Tv	�T����{�*��1/��������Cw���qɛ�A^si�D{�����ĺUw��(��'P_�zl�wvGX5 ��N�	�0욷�Ֆ��%��S��#�9�.���y�a��ԃ�r��u']���\��_��B.m���<P���i�xG�1%啂��T�Kn��=��n8�m/��Ү#o����%��ܮ��������F��,�s�o/+�>����/6�Nr�[�4�j��d��J��|"*s1[O!�	<�p��N|^c���|qJJ~3Pn�"���|{���W�>�	�� �IA���-��o�����7ӽ�dg�;��x�7ǳI6�ְ������G/t�ڬ���? ��ؠ��Mع��I�ؑ[[VS������5$�[��h��u%cn��=�+y���D�e��Ӆ�i�rB=a�8'�����DcC`g����?}n\�N�/�S���nw����S�����f
f�/d�]�Q���9a��8k~�5�����8�qiiY�����zztU�>���r2�x�T|cK�sA�܂Cu��Z��ʜ�.��:yeq1|��X�s�y�f�B,�*�/xTTTt݂4ؼqf�����aݖ�{C�T}� 1Ϫ�zt����2{ɠ�����>�e����Pp:u��0�1?;<l��!��6��L��.C]��'�7�k@�Z��z�M���vN»▄���ƃ'n�{c�K+���3��T^����Ymfk;l4���2IK:���Z�F���y���ύp�`�	�ps��ԥ%�]
s]��=��Y��Q�K�H���kii)�J����u��������e�e<�|cC҈����}d��ٳ�ڟ�N��7s�J*��J�JeZf����K������Ӧ�4�������KO�; Ȥ��8��+���[��OM����1d��[ތ�s�Z9zi��f��'N86H��av����{|�X>?'D�؇�g��z�P4��';�^�JL�w6d.?~K4@)a������/�`��,��	5��}�
�9�E�Y&���z"=DB�q�ev
���W�wŬ�y�Vf�M��o���;��4_��x��4#�6������j �3����7�p;�
�dM��V�=�����F���3;<��@���X�N��3����x�r.�	�"�j��WS7H������Z���>�[Z�L��=��~g���y�XDi:F��+U���l��纍��ɦRxT�M�#.c_��e:�S���AV]�P�V��]�r��~x�%EWD�qaa�e��>Q5�$�}�Z��<�?������8=$�����S�C��ts@+%�〖�&ݽ�"�KK��q�=�KA�����J�2�Z�ޑ�l��g^�n�mh���4�����q����Ǹn�&	C>��ի��Qi�k�IIIi�E3�*M����L+��5$���_�vU���k���zA���ck�|��h`U�0�m����fl�]�m߿;�C'˥����𷨩��b����#Lq5~�ܭ����2K!\�y͎1k�W_ÈY�~���V[KK���F�c�;cccG���_#V�Ha�n-	e��yכw�����zA,��b�:�V"ݖq�ۻDu����ļNK�Â��BJ�w�5�M���c��Y[sm5�ܾ����Y�[̯/�gX-*	=S��k5L�ŹС��5�ѩ�/����G:PU��eUB�f�^�5�R�M�"p�콋x"Č�s��f�8/XJ�[_��&Vc���	x�<bF��H��i\D��0�9p3���35�o\�κh�b	�h�>�x���Bh���b�22X|+�8��Bv�UO%�gM/��;|n�\��x�*1�[rFFK[[[�I)*I�y��*�����/0�M!=olq�|RaN��v(u02������ �N	z��>���엓�佦�������|��N�<�P������?}:�
�~nf2�����:��i�Hmt~��������k���o�ߠWh�qWO.}�hM��ː���h�p��ɞ�Q1㒢��ؚ',HҮSixZ��J 0Ay�`����W#�(ZM�t#Gj�4H�8Y�~�k�F����������F�'�8J�o%VJٴ5��#ص�X
��u�#6�ZJE��+>o|�}wu�hoM�p1����?�sƉ���W���7uu����3RR6�bb��|���F��H v>Gj�����
z6)m�~��ُ�	��Q�� ��I�f���y@�	?���0K�5X@�@aC�Axtc2N�y�{���Q����K ��B2��Nr�CCC�x�m�}z�;w���rw�P�(���#B�mm���W㫿@��~�Ğs�a?'7�vpp0����Q#<&���&b�i�S���_!�	���)o ����ߎ��G䈾c��,�I^5R�F����@�Z����)2K���՛�7��s���z�,� ���<��۪ �"7��W��0�Ar$��]��I^��{�C�s^�2ؚ�/���1��(��|�jg���}xn� B�Ϳ���]�B����Z|w|RxD�� ��Sa;z�^��8��E���|�Iȑ��/ �9��]��!� ��>�Yzy�z�\B�#��z�M�rvO��I]S��1+[�L���fϿđ-T$�����Y�� Ω���c#ȱ�c�{M����p
��:�����c�q�y��O�^�ih��MM w� F��E�&m"�n��o�MMM�ڶm[5�IMMM�W�\yB �����oNwJ�tP�rY%^��q�l�MN��^�b�;}��qr�]���y�8@�%�-�6�ܣG�1��h�c�4���ȳsTe=*y��� y/ Ȇ�S��NȒ�₧O�8�"��_�� 0��(�H�B����N#�וؤ�o���5��["�a�����zO�X�آx奄'�����uP��KֈO����N��{\��&���L4%p褰F\�r!We�ٗ-\\��&�@���V�?���?a���@�C�ù�7�%�)�
O����5׉���#O�43s��@���l<T�"�5������<Zz;26�]�0*�w�7��rԓ(�v�*+�탦	qY��.dGӱ��	uJ	'������� �!V����Ɣ����)6���c�(��m輰�)����zAWCpds����;�1ʤ��4�䎂�\�������p6��r|8�����oB�u�4�c��B�mY%�[p��98B�)ז�-����G�1>P�f�h"�ȧ��_-���bˈ?�p^��al49T8,�����#7-6ش�=vx/���e�m���䭚���vj���+�{!��˰����)�)Wa��\z({b�_�yv
�H��$]�l��i�0���Drd��F~��&�.�����̃f�ɕ��ϟ�5d�`�J�;��?��ڴ���
={z_tt4�����gyEk�����P{a0I���]
�fV�d*]B������V}C��c8� ����y ��<��e�_�v2���w��B����]뒒��A_O���´R����
��.��W�^� �zFQQ!G//�4f�.b^u�&]5�����>��n�>A�{�D3��7�Ƹ@�/A��du����u#|p箄zrS^OG�3�5eݾE�83 �f�	"�oA3 %���#�8z&p�4�5Cj��v�$�UUU[X�)��s㭶��K�kRF�
ڃhF�����5����=��ҕ��n1�v��0���PŲ(�И�����.�������'h�M}�c3(��|R6��@v�^��:9:x��L���`�
������ν��R���X�&9LL\Aa]��'Y�JāL���������
�|�T����T����P�[P0��hIE�Y�N��<G�ʠ��̸��QQ�A��ܾ�*�jhԥ`�F�� �`o�����N������%W��cIE8w$�q���� 4�����Q%m���kD[C����������&���?�:9�t��9]-V�S���O���эI%sk����)�{i��Wިg�kHf�A|���� o%�r��9H�8"��f(�nb��s|N��aTjyv4���b�I{7���ĩ]�=���Ψ|���Ƞ��B#4S!f[�����lH5.������^����0��ٞ��M����G]jG�ۓ	�a܊�X�!�|����ݲ����4���v������JI�������5p#|�_��y���Yǃ�W����Dk�@}{��}KK�1�J�y�N�#E����Qz�ƌ�{��馶��V�Em��=_� OC�NP�7���M ��KJNEEV7|P9X��G�N�#BY��p�c��!����T�;i���v�S�pW]]]���ӯSɧ_*գ��^GK	�tJ����K�.5'��sAy�;��K\��Hb��'���^�Fxꭋ�����A�˗a�(!�f�)ih����x�Ǿ��o�Aߚ���@��G.=+쯡0���ЉM7Y>���Q��o��Aà���3��#��W��[��	'�jio7t��K$�"#���B�蠭*�A��y�tP�
ı�pC����@��<����6��@���ḥ��Ī'{w+�7"�_��O�"��A�l��^@��KӴR�j+|�"����s	��H�������w�`�ñ���'O�	��d�:��2���dQ��_�P ��J��E����QQA����Q��_i;�;�������8���0�p�22b'��*~�Fm�7�����O!ި�C��r��`���OI��
�]X�ϖ�\�?���������
O��Q��1��Gy��-|s���|�'ළ�}�?��d���Nk��4u�Ij�"�j�˪��n%Y�D�.=�]��;��������,�߅\�b��RUQ�v�À ��,�έ�*Z��J��]��c4�s��~wwi���1�܍��/�-��O��Tg�����r�f�M*U�ژX��#[�U��Wtm Y"��ȑV�1G���:��p5KԼ�}�v�g����c�z��o���O��wUB�x���=��qqqe�9z���F˱�R��Ցk��][���a�6( ��Z�Ƌ���E�a����dq�΢��Q8�ic
������p3%�`C�cN���&����y	��[�C�f��Y#B��,���+��xW�����������/q;�>:r�%υ$�-�p���hڪ�.�)���|�U�~�t�˨�ïtD�۾���s��D/����m&^*r������W�ᠳ3���,Fà3S�c�]�Q�6�K�OÚ�zU��r��"|��^N�N��J��Z��v�'GO��`�V�RC�<�|�͠��[�F��³�,HO��'�QqD���S�Rô�N��5WA�:��@�섟�c$�F�������>~k����^̐��-�G+4�_��{�I�^VV��dXGR�*��3�'���W�[�E��0K=���o������u��"�#<�P����%�$���9j���8�\�)�9@���/�p?�l���:|��2���zmz{��d��8��!�k�,+!�d�x����h�@���ts��Ç�e?�5��.JHI�N]'��]ҧ3�
��U|)��Zr%̛�ؠx�r���y�Op�g
v����-װ�j�R�E��z;;;��x�C��4��>���<>*k,�wVhn����ts�������:�#��~&;�k܊��+l��ۖ=5E����%�8d���z��o(�(#�af�O��\�#�W&n`0�˂H��'C���9�,u���Ӗ��K�76�[��nl�&̍o�!ͪ���D<�=@9%���X�c��Y�_���O
�d�{���1��%c�Nt�����s���3��]Z�0%�	�[k���ց݆BW�z
>K�/ �t;#8����g0�/��`\Hو�Ʉ���\H�d��:9�GguÓ{z{�е*8��,-�G����*�w9xm[�UZL�d�0M���XW����k/�}|�9v���wEk�줋�ǆ�[X�����M8D�~�h2f������,/..��/��Cl��XX��*u�5�u�[�������3�!D$�{�"��Ý�h8%�ړ��r��s��
k��a	�!>����5��]v��_���(SN��.H�=$����?-
,��0ӭ]����S��ٵG����h�*�8��u����"��r65%���n���U,lޘе�ʝ|ŎP�&1��V,���)�G���E��k�ЉOn��|��^<(%E%5�@�9�l ���6��bI$} V5�Y��qgF�������0d"&�n`�s��Y�x"�p�s�b��;����E���K���b>o *��W`㊮ ������%�'�z�9�O�[�����v�ݼ�vd�Xb!�ۋ)Oe�'��v׸���	�Q�>��d�iral���V�������ct��g�ȋ�}�PGl�E��MI�9��'��o*ң��x+vv{,Xʐ�a��g������X5���^,�>yD漂	� ��t��b�x�Y�5n����v��&af�E�����y��m~� ]-�ޅ����<��w�L7�Sh�3�����ĆX,P���J�T��R,w;�Oc�'���ɠ��q_� ~vn=H׫�I��酦�;4�p���R(�ER؜: ��֍��&ڟ���bF�Яu�t6�Fy� ��>�����
�VDB$��b�����B��d�+'n�P~����Ǣ�֔c��K뱛���Ő�-	�'e8$ T�����"3I�<������s+��m�ӳѺ��a��`3�TZ�F�B�R�,|'((��y�/�
� KG�����Q��!��t�7YF&t3
>����
��TCfCB��K���)����3)���Z��v�H,O�A&ka��czB:e>��c�~Ze`Z�nߧk2�Q���V��{��ʎ_�;~���-Jm�+e��%��_�hZy�aw��/L'�f��m��][�s<~c�"�A������c��Z��^�y���Z��]�v�`����2�d�F:(JKǪ+�U�-���k&cnL�sn4~^*2�<�B2wN�(Ȯ({z'��[˄�Ol���E�uY�*��ܷ��`��; �^aw�('�*2�6(J��P�{j��=Y��׶K�T	��\̨�yP��"���0�	,L�0��A6���P�n���%�k���J�'����u��p����k`�ƛ�z֭��T,���C9�� a�-��jXX�ɡu��������9?��#g������C[�������'E&�N�����|:��zn���'�`y���1.�i_1�P���G铴�ie�{����ͱ�@;x�"��`�!Nl�9�}8��~�F5N����`(_���-��Q*�n�*~��Pd��n�I�4�j���N��N4�\��u}��[`z�'�˺м��ƚ�i�SLr1�r�=e^,��8�;�*�e��M^O�x��˓���L&���e)��s�����Ċ�z����>�#���nxF����qUBk�-��[wͼ���B�݃�i�2q�W�����B�a����(�ޫ��.��w {<�󯀖9j�~��C47�㡧�CK�65@�ͣX��`wHu����n�;&2XC���߅���JDkx*LW��^��Y2�����  �b"|`��M|���V� I����m!�w�ܙж�~kN]�R���B1�ə�aW��ħ��!{*��������n�����q�"ڶd��`��7�����0P�&L��2=w�䚌`�ͬ]w}}}9�t��B��z[�Ggx�����rH���챪�[L%]��~��c�\B�a��ݤ��g�}�HUi�/_ᛛ����!pMd��&v�BvP���� Õe#�X���G��qn/���#��� �����W�9;�̽��f�S�A�&O�3�˄��DH#C��i6��򹒯�)9�Z0��K��ȒB��V+��\j�ݸu�Փ�?O��=��%h�Q'C���E�̍Aڂ�n�,C�R���-��{��Xab��v�<�/�{���#O�6�-.�D[oW��=;6:q|,�6ۛnT<��L �J���={���ңpIC7<��~ya�F��Зb'PM��g�+�U/x��﹦�(�A�aѹ�,#�p1{��R�xZ����ʮ���`pa7N&��?Lv�|�> X P�]�ש�e�l�Z�}_a��� ��!�\��\Ú�3F��.��F�v]�ip�u�!�����t��nd������q��R�S!H���3���{�����8��&�l�\qx���r)�q��DF�چ��A珮���û�K��O�;�o!ţ��$oʨ�$>���7�YR�}����
ѷ��� ٥=]B%8r ���I�,��2��رKHz!��oR��}��@>|L7�/��=��%�J���>�{��ڱ�島�.޻�
�U1q˨����6]����9U�8y����qcK�0�bǈ�,�co�{����xC(L�P`&�#�Τ���v7�y��WQ�o��/WM��jl͝gEK�N���v���pQ^m��'�K�YnȜ܎��S?�+��?�s�E/pi�$ab���Z�7�ї�<u(C&J��[s�rKmv��&�1����,�aDb��'����9g�zۮ�VI)����~�?v2��ӺR��A�V�0��Rz^�nfk��J�$~E��/d�ކ_;���,Zs�k�l�<ޮ<�V `�B�kW���l�&k��Q71���{��u�jۈL}Ux�Wr���X����T2mJ���4T�Ԕ/���z��B��U�3/g/�kV���`<�g�� {��Sj1�Q��%罔Ґ!scX�W+����<���F4�R��RR�����{~{��|�~~���>��є��E�!��C�j�x퐏/ݤ�������Lf��L���m���X���Y2��E;;�o�ꬃ"��ܾ7V��ڟ��م�4�D�ѐ}���S*	dF�P�q ,��$��ŋ3���c��Y5�-R=�Xl�����V�o]���+�l�]�B�5<�e�Q4�
�f��[	KX.�/
���eI�B���(���P�'�"+��.B" T�bz��^rE�e`��=CDU�h�0ǃ�F���aU�*c��At�7�ևi�b�-!U�w��Xg�i_xd��T����{���,�/H�Q�ɠ[�Փ�z��Y�E��a"p���W�An������?���c�E-�.6�B>��I�pE��VV��@�=8�P���)� ��kY�
�@�rz9֛���B�$�Uf'K���T	��"J�ޥ����}�O!�� ;�b8�
�*�m�A��M�#!��Ȳu���T��+;��e�@������_ L��µ�Bڦu�T�R����s�� /�r͡�N��6Q='�u~XQ�����
+�&�j�B�4�?��Ȁ	1"�(9�PA�T�!��ν��4ϱ/�h�:��ѹ?��c�o�����E{!������-v��Li��MW��rB�0��u�>(���.h{#]�K�+����;�wuD`����E}2sEk� �,��ߚ�گg�"� 3����]&X�T��G�#3�N�Q&�E&úU��@�����E@g���#�Q�/���N�)�����K�ݯ6zd���8��uT�(2l�ձ�ETok��(Ah��x8����Tg�|Bi�@�܃���RRj%�F��l
�LI����-*�����S����׼hR2:�p����\B��
})�-Q5�	-v{������D�jb1�x��@�j�U�$ZD�kAFYꉄ?}������i�R�m�SG
$���_�m�F�L��2f㱵�k�s?o9��M�"O����,DkM�կ͞��P����&�*cn._���<G��\��c�<�E�<!�I�nIMM��D0�<���Q�h�/7g/���Y�+̣��A8�������� ��0(�z0h��%��s���;��ɒaø�{l�C���=N#:���d���'��̴Q`�Ɣ�@LI˜�Vf<Y�-I}�S+A�Vgy�'��*8rc�Ҹ��}(�^�-ND^pشdk���Κo�?X��{e�]�v��]��s�[��7 ��s�a:��Km�3��D��M��g��G���eB>�a��n��<4�;�4û'����N�Ů0�#��b$�R��c:��zU}���6����]&��{�����Q�g�*�G��t.ݒ�_@�Cz9�TjFR(`��y��@�Co� ��y�q[r�0W�٤��E(� ��Bor-O��@OG`p?\*�͗��t��ڄ�����^K0�-~u~�&@b݃����H����0m#ݥ# ��Ijcd���vy��Nl�XS�~ '�vF:
��Nё)�
M":�u�[7�x{#��ח��d{(5"�;j�uCk��j�A,F5�DÖ!8�uk/���]y�))�"����XE��))S.�IX(��'S�ڸs���9���8��$��b.p_���71�o�ޢ]%ɔ�/g9�q㑰���t��F�}݈��j��	{7����<�=��6�vԙ�a/�W4��9�,p6;F��,�NY�L��C�H"�10�gv��Ú�yO49��8���W ��A�1A(( NOBuP�����1����?��1�v#Je�<��GO�B��i :����sB'�2|⍫����GE{)	���$�8�}(p��%�#Sc�
(r�ؽ�#w�E���4Me��
�Η�A�2����mB��!l�aaЂ ���,���3�9<��:��C_�f���`7�\2�RRp��O���޽Ϟ�>�Mݣ4��� "\O�B�9pO�k���^3��.B���M��$=�u,��hc��I���K�J]J��:� �މ�Ԏ�[�J�ch�H:lV������}[ی�v���A���0�ފ�X�� SJ�	�_�2SR
xM�A©�f�	�j��=�Qs�4��E�0~g�&��՜�;9g�L��EŚa��;�Y2cA� vږ���k���,��:c-�*T��^,�0�"���ee�+6G��s�5'�k,�x6�f-R�&/x����~�s�>� 5q�����@��X��Kg�B�U2�5r��۳̀�t ������ބ6�̧���@v�9��-4^,h�����Z�E���uFL�Jh�C�7%C�L �P�!��f��6D�B�@���|�w��*u��olđw��uM���9��"Jr���[s@��A��f�u�ģ햋X����7/L��#��t���PJ#-������Pv#���h��b�M.�T���If����9΀�KU"��<R�5�2_����W���P���U��$���e��A�i���~�ͬ���	�̿At�g�vE��sT7��0�J2�g@���}6B�P{{�:%����х� ���Ċg[�%��(̾�rU�"op%+��-Q��n��* ��틸R��1!�ъe���u�5�]�$daiQJ�T9o�嶍#7��3fDjf.�����P��)��x�&G˪�����	UHf��[�ѭ�X*/��)��U�"/
�1��t�zz
j����<1)��lX��"�}_���}8Fz�h�S{>Ta�����fe}�@�O#Q[��ezή5ǜ�n�[�B]�P�2��|��xb�r����/�M�TP���Ix�m>�����j��<�-�2К*�"��J�וރBp��9'û���U�����s֯S���'>vY.�S��U-�K�F�����Pl֧6^�~Nv&��@���*� �G%��{y�>A+���i DT�F�����Ŋ�s�Bch��.6E�1�l��{�ӧH����&��:��B�e��9T��í�|�ڨ�0�$i��:l�k�Y�o#J����Ek�����b�B��:����_�]h�X�y����@�g�Ȃ���ݪHSl���r�e B��nrx�4�-�3H�B��]��HI��慺6/��+e��łJ����2�f"��@�+�T�����N�-����v���O �:��-��}�j�3�������AJ���	�h��$^O�h!)��>#� y��+�Q=�ѧ"(q=�[��k2{��	�Їӭ[��n�ГAbx�	b8 �d_,9>8\s��ğ+�px8<]�^p�93�!�W`>P�򂦎Z���\�(�l׿ї�T#voDy>s A�Q���,�t����h�a��&P�E99�|6
Xb�����XI���ahF����@� �5��.u�FyU�$��jbà�7�$.�{Np|��LFX�ٶ�|�B��V��A�G����wxRJ�X���GM"�����r�r�?6�bM��tI")\��޽��ӈ�h1��R�T Ha��ޘ3�͍t�DK��ܱŔ���R��H�G��[2��<����yM��m�6�[z�B�߀-���#���W�h^�o&��}Ȏ,������q;.f��q�� ��RR����޸�R��PIU�Rk�YpǸ*��.�����7f�1c�h�}����	1P�11_QfWd�Z	P\����m���N���q��Ե�ի���ߖ1ӝ�擲�D�KG	��@J�[(�<�J�Ғ#�8��/�Z�f�@g*�j���`��S�iG�q���z�������s��j_1��:�CS%���ja���T|u<8\@ɼ�a�y?��M�%DG��L�_������N��Z"�&_��'L~��F�H|ˢ2�xwi[�W��p�_(���aY���w��Q&��ZT'�{[������Q(j���k�������L'�b�h�ƴ�4�ˍc�4[Z��#ɘ�����4�m�S�2G{��%��d�����"Cs��ڇ#8}z���LeJ�^�'iR	<�`xz��ׇ��mff|9T	s��k��D�7�f����ʶd�4<}�H��baK��\ZJ߈vK�.D�<.�Tnh ���3+�{v*E�%"�f箯��r��U�!(~�����":�()����9;�>Fr?߼0�8n��+��{�Q������� �[K$�ؐ�oAD��]�F�	�횃Tx��X`|�6R��'����4��bv��4 ��O����z~j�ō�A�U7̝D���ǿ�datLdr�G��k����)@0\#9���$z���ȉ����KԀ�/P)4� �K�K�d�����w�y������*ꤦ|�D3KJIф\SD7���-���I�d[O�PAUu�Fy΃-,$���1t�[�r���XE���Đ3�m+)�ǐ�\�C�^����@%��d���(�aX8��Y���yDKa�y1�⿹B�&�b��W����A���G!�� Q��B��L�Њ��#g�=�u���ۈ�3K(cÏa�d�g��$�	�;*�\F�LV�:0rj�O/O��Ff�w���&��U1/H.��qr���Nl뱡{��q�oJ��i(�@�J�|⍠����O41��v�f��e <�P�n�I��pBV�D�#j
Zxb�W��@U�B)J�fba0�XJJ�o'^�DB@��P@�̡���������?��ڼ�ī�H��}iD--BH�kt�5�x�K6�T�n8��r��F��F��3�-J�) `���ū���c�"M�j�Ry0�8hi)"pE@��!{k���/C�ՠH z�ӆ��Ow��5�g��l��Ql���1�)y4o�_`��|�B)���;�Ġ��Ea%~���0Ū\�:=E|'�'��P־|>h0<b�t!n��<��n��%��k�~�
۩m��aK�����ܡ��	"��������b�w����k �O��JZ=���-�Q�3,x����\fU��R��%�]�-��ù|�Ы�gx��e]G��aySD
�Z�>�yM���P����}�d�úsPH*"��&O��z�l͓���+Nq�{�\1��)'��_L��=�ɞ}�����V��Ő퟿"���T�SY� R��Bp�a�}��	��AaXR�Z��y{���"���c�D9`��N������tþg�#f��o��RgO-�1�NhLkN���6r> N��qWP�����X��b�����XX�^[�Q:�B:bhI�҄�t�(��#��w�?@\M�nr7���>v�!T�A>�.�k��m�4{^,�c�� �?�AJ	�����BZ ��dJ��&p�W����R�c���6�2?�H �H�)
��
���jQ��XzF����M���V��c�T	��(�P��S1/��+���V�S,�(A�{*�p���Dk�EQ�?B�C�,D��GLiV��^�i��A6�ҡ<A9er�J;1��j#��E�Ƃ�.���!�颦2���3�[|�d��=5��{�Q>�����n[S�^��tA��^�!,f7J�����K�W݀N���X`���Zrü<6[c(h����Dx��(X��%J���&��f�5�l5'rf]����it�i���!��1=T��]ʓ��QL��.���rSj��]�Ҏ�Rw��J�Ȃt���s�ʮU��s^�J�ɡ�����k�x�)�J|��Mtf;��b�E�ޙG9|a��Hp9��̮4=%r^�5g^M�K�$L�	���ל[�����\��%:� -.��%z
������e#d��E�����܌r�5-:@�7�Μ�G�&~�76��R�0�Yy`�M]����\)WVn�]�<��_t�~}�.�j���̶�α����U6I\t�ٰ�@4�/2�Kп�Rb�Z�7F�7lw�8k�3����z�����~�9_;����,�w^ ��m._��I�P"p(���3v}����{��p1{Hمr�RB�7a�'U�y�乙d1�g����M�ްz�w����hhTR�2Q�=��w�J�M���1=;���Gل��T�R�JN,�h9����I���va�6�'�#�؄�~��k2��ƶi+�	a��J�h�f��Ϝy'���5�XC�X���2�f}?�N�k�F�ܓ�_I��N����u$(���ޙ���m�w?i���1�I�Y�
�R�[C��0��ӓ-����~q�����fʦ�Q�����,�;*�/�h�{>�����a��KB�oUa��9���:�O��f�3�_<Du�������ϸ��|�U�k��$�;%�z�~
�)ﲦ�m�f�="/$�\;�y��>x[��5i��b�x#�҈mG�{�'� Q��}Q��DW0}�~NiQ[����oJ�s�)�?ij�A<���%��B����.Vi%��Rz�Vq+nr�9�s2ւ���M�
?�0� ��<je݌�$���0S��ɏ�D�����<B��-Mw~���O��]�J�_�F~�_��[���[��[�i.\�W��w��m�.XDQ�q�[y�H�j2 ̛����Ckm���X�b�:��I}iz���Cfˤe;A��or�c�f��[]uߵ�L��g��V�~�]�f��=>J�̇���W�g��j![,��%a��o�����뉕t���Vr)=���1�1<ہ���V�AF�;W�u�'ӹ�@��:p�*��4��;���ۤ�9�T��,����g�Q�{h�!��ε�;L��6r�
N>Q�~"x�r+����H"JYb�Ȥ��"�������hh�ۄ���-Ӭ.^X��7I�d}߲L8��8���������)p�9>=[��.d��UEe2/��������?S��f�m��0�zb�t�~�����؅^��Hp[�9�����\���T٭D�IѾ�%��ғH�4U��]��E�$��$�$�r��땢ͳi�<�\&˰%���V�%��.�;�%��z�D�(͸ub�7��J��O��ʡ�>
�����z��n"���F�OYm���qZ�Ή5�-�άƄ�X�k#��ȘQ��5\"D~��:�}�XJv�d4c2�&�ˈ���W�d�*¸?C�������7����`Qݜ�$�;�Efx�6,ʝ�$�o��b	�#���]Xk����S�"?c#d�~����E��lլM�p�O�ƣwF'l�tRQO���B���½�w�p�!�u�c�O1�a�CG����Y�ad-`��գ��DV��"���D8*�(5��5����b`�f_�[x�N譄ӎ@ �W���/kV�m's�f�b�0�9&�-������#)�S25��I����\�.U|jIg�����s(S�����\�b�P�	��i8�z�^��T���{��2�M��\\/�0��h�Á^�e�w~��r��4[j��=�8�Heb�ף3�	�G�,�Z����6�,)H�N*��3����?[+�"R<^I��d �(����*�����:��b#`8��⩋B��a�p��)��h�Pb(���D ��؀�Cirb�Q��g�=�2D=rt��k���#���h�Ϣ(����a���ZVc^�lO��Y^@�D\_�����?��̦d����2,V}`^������tl��JG_},8������l�p�A�Z����Tw���I��`˻�)���֬N8��5�L|�k` ������#�qwҲ���2LC��ېc��X�	�C���74���^��<A�Epwܖ��� -��J�5g7,^��I_Dq�X,���'��*�S�>(YX#�!��˧���'�7T`@���ԍ1���!�K��*ޤ9Pg7k9��I�h"O��  >Xߪ�d��ѝ�E{��t�oM���=����͘'5����	�*P�:ݠ*�Ҿ+Ӿ������у>���42����X6#[r�=��܉��zS���/醢�PP���砲�i=m�T ���^��y���f�_(�}�I���
�ӫC&���_�1G���w�7D���Q( 2�^��� 'Ǒ��"��-b�M_b-��'>0��h{��e���&��w��#�n�6�<Z������UNa�t�ee��}Q�T}�̽����/w[�gK�R:�R:��6�q����D�����]�8d.�Ec��R�葄C���μ�
IN/�`�9<��`Mw��w��"����M�*'�
��8�m��?�l�#��Y�N����	isB��4�g?s�vH�)� ���Mɇ��w.�����s�H��-I���PZ���q�<�N��K�͠}@o��v��)�"�KϪ$� ��[HeS��b弦����=s�7
��Џ��ӲeC����>y����2��TQt�Џ����x�DVq�V���&������1mM�yх�7uIs�^pb�6%�.�w��b�_���5��ˇ���ks�c��0<�`�������zJ�K�P_���ғV֣ϖ
ΜE�_���#1�]��V��hY�װrm����������d�;i�*�̠ٜ�Z���FSk�o�Y�,�E��i�P�saY�3)��#�5�#^����p�]v�G�x��@X�+z,�E�b8ڽ����k�U�u��L=>�����M�@|�S1{�'��K�>�PZc�_o�����0�w=�����#*}g�� !z�[����m�洠�E� �C���"�i��C)�м[m��כ�V��E�
�)��a�䂇�	1��?δ31o��cV�W��t��>7=�˩Aˉ�Ik,�I��{�I=L6���	q4@[:�>��&�ݦ$w�#S\u`���L^���^`VG���i�E�{=���ށgk�(��n��_9R�Y|ta�K3b�(��2-Z��\����#V��"�����2����RP�d�	�ю��b�W��:7�cRЌ�AF��V�[�C:�?��@W�#�U��s<�'���_vOJa�W�z�����R-�w;U�|�R����
����+�2���	��
�t�c.?&R���*"e�u����E=G�(ׅ���Y�����P͎�&�T'9w��awH"9�����J�ag���1)��`=��b���`��Mj���j�䏢7�c�{TF�t�ؕ*���+81!ăH4�|�%S/��������g���`�M�c1t����=1�Z]�J�m�E��ߤW��`�0>t�&T�d��Af�&Ν���]��a���q=��7Zf�d�AN�t���B�o�:��?�X�D%�%��:����S���g�,�X����#w'�Vj�1-IL$��6A��������� j�&ws��9���W�3f[���T�:��0Q~)@~�͡o�Q�>�E>��|�7��yơ��(�؞k\?q�G��
4n+�B��`�u�"~k��2��=�f�����?~:W�׏�Q�h���%�a08�����.�W�ὶ��7k��>+�t�����X��}��O%��2�r�I7~�N�O����n� ;}��l�S���k����s%��9zT�2�<m?��!)�u�������wI뮂��ڴ1m���}R��г�-F�"^S咨�Q �X�� 
�(@�-�����Ǣ��f�i��齄�d[1��庣ia{�FX�����=k$�pjf����A�a$�0|��""�B (Ķ����Q��,�Pb�?2��)���-���tP�^��&��<8���]��A��5Uts���tG�L��v{"4��{».�����׿�`Q��U0ڿ��-��}·5ҷ�J�Yq%,��`�G��cR�7�8�L�u�b��=<w��?������y7�}��Ӳ�,,���Do\jf�fj������L���7(�u�!��.l�ݚq��2��XƳ�d�8�{v�H\3��O��n�%�9�%\	�ɪ+�L�C����m&������E@��*uT�FS���p�2�x�)��$aV��]2OZ�k��Do��e^�#� ���=�a�0�x�=l�JZ��т7z|�C�sCF���L�/Y(ȫ��wܜ�]\�����/��K�"�m} ���4����?��ݒ�iYJZv[/uX�4��q�d���)�C��W֗m'��!�60f���y���,�9�u�x���P"썰L�s<v�-~���W]�{�Qt\��{� ��W��}+���6��Yf�%oN��C�8�	�id}ѩ�|��Mq����~��R�� _���1�O��"� F�lP>��P�K���UH����4�{V\�%�2�/[;凵��_Hާ�}���W�^<�G�����iO\3�:�i֓*_�hį*�y!gxs�2��iECa�GC��8�������y��Ө����~���S�%F����ע�zCsZ��l�[.J��K
���7�e�.A9X>`��1߃=$_�(/_�jݐ�鈱��2��.J��_�����x�����{S7ѽ����ݨ&K��n]*��U#�ܡT�d}ZdK�Ie)B2b�F���${��[��{�3K�������}�ky����9����u��R1�Y�ʪ�.��$:���}f"�,TƗ۬��#�9-?X�ً�o���S�ş���q&���t���P�{W>]x�25�����Oz��AYP(:N���h/x�$z` ���q�� <��??��� ��h�|Q�XV�I%���)?�(V��	�_��\�ĬF��g���aF&9�|n�������0n�~L8n�(�sUvu���P d����4�B�8MQ���v�v\�ol���[�;��D=�s�`���\܏Tt@����}	��,�|g���2F��q!�����'>L���v����TV�3�ƶCd��C����?�3D��%k�Ь�2-��;Pg��u��H�1�Ч��eʔ�U�언�1�m2,���pzɇµq������:�8������߼�i�A�[�"��Ҫ�f�	S�f�q$�+��xm���g*�z��v{o��n��|�_^=��;%,��(�J�A-��7,����)Ѵ���V�zAƈ�����X�U4���a�{�[���ŝ�l���h�%HA'Lx��M���p��%#���8ytY v�ջ����_�C'���c;�<h����vo��,���ogw�J�ݵ�s9�aK�%�����:>=�:���-�����Pʏ>qU�;���v�H�7�����r�[T+�e����0
����.�w��\�P���{]h {�wj�R�+b���8��^?xP/�������\�	�Z��oމG@H�N>g�yn+?e�6���IGcQ������ߏ~��b�8ˇx��(a�2�쁫x��n/�����~�7���g��������;�xIc&�(�j��5�عk�Լ[�e"l��3J-2�L��1�TlDT���@���&s�k�;�jZ�'�ۖo�#�$��#�AU���-��fN�tɔ�Gզz'!Q�����|��E�<2���]F�O�nq�4G�z,?����Q�)��C�;+2�=�]�����_4On#|¶rHn�s��<�S	��Tns��<��/�����e*�S*얃StK0o՚��M�y����v'�a�:��:Z��j�Ӈ2߾v^��2�1�4��?;�>�8�B+ϟ{F��	>�6�dՄ�����0!��~�[�H���6k[T���>Rg����?���fi�� ��a�Y�s;�~s{��Դ���/読���I+�������\W>R��.��6җ6�o�����t���hU-�����'ET֨�%^js��{3[�]�r����G!L�$�J7���fq����
o��������2�[Y�r��5|��~���'ܡk�@g/�Q�^��)�K�!�v��mxT��d#F/��a>�������ˠ{�!� l�r�@�IEFF"���K��/>�\�?�Af{�31
V�UQڣ�y���x�8�[
��q ���?����n�H��Y͟ϧ%0逾���1��X��8�!��rC*	~K�_�t��
�'�����\��g�&A[�@�ۇ>���`�F����]��k��`����֋h����!U/&8m�^�88Nw�p�=g)��EĞ䎛��1��{ǟ�=Ϩ��Ƕi ͡=���v�-�9�Y� _�:iL�Αr������f�8[Qt�G�
BԢG(�ooq�(�4�T��w���ř�JrV��页N��{��z%�6_cCuh� v��N�h�5������� ~T9(���ufF@0/*����F
�t��Cg��u/��Ƅ^�i+��]��̞�����w5g�����q{���n �_V�`���}���/{�C���K��j~'~�P�^�`p�	����}�J��x��hi1A���3~M��5�?j��8A�Q:������О#����3ɝw���*����e4�{����|YK�xf���ȂA�}��5Z�1�x�V�{�x�ۇv��E67�-�%����:[3���
j�_#37˖��e�A�^љc��+|���绅�7v%�Y)�H�]$��V\Y��;���"Έ�g��s�����.ϖ��*�f��:W�3tz�a3V�b��
[}'�7��~5��S��+��w�Q�z��L�Õ�:H��i���?���v||��l��v����3�W_�z&����+�܋����P�D(��Y6��1`O6�w݀�1rɺ�Z��33�=�M���WN� �Aɯ�w��{�r�$�n;�d�J �����\�Aܿ��n�7JH��jqlɯ��ۆ� x�qr�3�����4��,����Ƀ�3D�V�]626>~�g�n�oӳ����W0m��6��ݼvp���qr��[��ttt�<�Q(���5�y����8����3բ\KG�[�7�����{K�y?K^4�w�.J�r��vWa�%^�٭g�Nsw�q+����0�?{�`y���Q��MSS37�_��VC�d��Y6ZXZ^ o :v�hR��rf���������`�#��K��p]H�Dg
�:	0�g�~@O�o߮����F�p|LR�q++�����y�h)4�/���7�󍊈�TV�I��T)K���mE��K\Nh�G�`544��/	|�?F˟\�����<�
cŅ��w��޷�m��8,�:�TW���a�`�B�~󒕕7o���<�������^^l�nS�C^���o۶@E��}���	��U#��y�ɷo��z�*�T��ed��)����SYw!�A*���@*8�^8/wYp���}}g�A�&�']�2�!L�"��1�C���ʏG�C�y�ոp 8��}x��?�g�� �RR�{)z&jaGɖ� �l��߄��%��,�)��I��W��&�xOu��9X)ӌ?�zwo�9����oPZ�=�o����
W�kRbl8�~t�¨�1�>������k��;�	B�"��ޒuGS6_�)J��g�4F���8!2**%��7��0j��#4,l�^-�/χ�� %F���W�<Gg�j &�2(^�_��R-7DY�~�����ᖰ.���h<D;��U!l�0���q"��~��\��8��Q¨
��c���22^ەm�������c�-j�aP��nn��E-���p$�0�wPY%nL'�	��vZAf=��+%�}�OM���7��-��;x��Q����e~o���B�@XVm5�H��ZX 儷�zSB��x�!*�Ke �Ƿ)(�E�v��M�ܯЪRüL���r����8�{/hT�h9��'<�PSS�0� �Z����7�4l o����%^�G/Wb��74A:��^�y+-%u֎�S��;f�?��+GF��	����N�M�aPP��nѳ�C�po��R}�֘�ty�ѝ�B�ah�L����5R*~9�V}J��hSj?��kU��P�}aM� �DT{5mS�Ȧ_��+E$Mm��!Jlt��N�H!|�������w�⇄��)�� F�'�OP��i~���+G:::�jy���NKo���ĖE�f��`�_�V�+l�w�@��w?_o�GRP@����`�E�{�:�15~H���K��|��xzf#����'��֏�w�F�̈�LTd�9��AQ-Rm�kC�;��b�|�w;��Խh����,��M�E~���ٳ�P`��gS�~IY-bE*���.��Il���uhn�8W�cP&�lݺ��J��ᳳ����{��,--=	e�:�tqPP��c!EWl��o޼��f�A0���Ǧ1r�R�L��&�������?S�G��5�O� X��III�m��7Ç��9�}�`�S�������G��F����36ZW�\�����ڥNa0T�Er<���K^ꤲ�x:�k�[�q?G8���PQ@Dq�8#7w�xT�$?�mVAT�8�E@T�����C��^�z���mTW�`�!bbb(���AHnÿ�A]q=4tP��U�tt�6��dI�Pₕ�Xq��u�c�LR�Keu�<��Hz���=��H�MBB��:��?&��Y8�aF$�V���ݻ�#���75uu�4�/��j�݆e��V�ɯ]��!A�9���W�� xm��~XI
�J�8�� l��^�Qȉ��[=������Nԯ�N��:�E]�h�����Ne�^	�f�?v.٤��o������&�w�6��wM���;�ĨYH���� �c��V�bT�`����	�O�IYs��v
Ӫ*./Gإ��p�֬��3=�/�~�/xxd��}��@@��"�1�i�U�����6��#�;65��3�Z8�kC�C��H�̤�9*p�~�7!׹�X���3��;9$Ե�g!�B~�RL\<��8�Lޜ��Vܯ��oq�M Pn�|+� ��1�o-�J��/j�r��v��A'� �)P,�Z���QN�-=��
(�K�@�v���6�_��|8�����0�.��z�O�����z9y���D �08~j�?BN��eee�)�I{!!��P�c�6_p$=jw�zwJe� ۉ�UV�$$nhۃ0���
4p�d��&���1���y�%��)����$��V��0)(ꔛ"� ���0����y��ֱ;w��C�W1������]��!�\B�?�DK�cP_�q8JF��0��&<�(s�A	H�����qU��2<{��'%%%�C�_�2�5�΃���Nw��f��]��Cm/�[�(��7���9�ԴV�|��^؈b'J<B �nX@�hn>^߸��A�����4�h�O�}=:�ޕ�O�qm��O���=b7������u�ʃ�B�O���_�X�*���oGFΓ��v��(P�QYU�?8����l�j�%��u!�7��x�-�G��B��נ���~����Є�/a��j�yf&�zoG�.%��6�Z�2�[E&i5ȹA�C���e�q�"��t�]��\~����PW�'#�?
�h�F��+M����=��B���0�L-`m�av>`�p�������^kQH���$�777\j�;�����88�Z4�K"��D�Q�����jh������+�H����;��	tĀ�Jf��k֤�:�w���³�S*Q���B�=x����I����޵��TeX��_DDD|�"��	"(�6k�k�[9��9�1�>=��kzzZ��1��Z�I��O�I?x�g?>'~����I�T�L:�i�-��x �s���>��m�"�4���yV	�P�u��8��1rLt��U.xY_��}:"�N��]�Gq��~�<66V7T?�6?����h�Z�@�;�cǶ���,Nh���`��	
���W;�;�f3�>�����5�-b�#��+�Fb���¥��Qul�I�C�RS,-,�n~[�8�ڝ�6`��|owE^�(qd��y1(z=	�P��[����]�%�}PQ���/�J�px�&�Cx<FNJO���e/�|9(SB,����g]g�D �6��aq0r85� Mb��e����t�;d��}�y4f#^������C��%������]�=�3 �ǈP���t�@���եIe�!��a;3oUH�u�j�,x���tq�sL��:v�^��+;�I�j�Jص]�[ߛ�!]X�{���?d�l �==bY������Z��^T��Di7~�X̫{$��AG:+I��P� z��Q���p\��ʊ���
���#4^[�pwH���e��8���O�M���������]:N��{�.9�i�D��ދ^�qT�$~��Uww�8�S�(������f��P{�vv�FG,��A���������rx�}"�,��-@X����1P��޵,��E��__��9�D��r�aEu�c���GL�ʬ���I�A
Vy��9�x�}��ʪ%�t�?�B�MM���kl	>�� �pB��~�Y��8~i7�&m�����6�jj������Ux��9кT��E�����Y�?qb<\Z6W6��_'�%�իW/W����l�����-�L���n�@uxF�[��:i���q�C_�cVfݥxF	"��S��੿v����v��jDQ໫���÷�Z�lװu?I�@��[�'��K��D�|n�6�������|�<+1W�l���f8�Z�����靐�������W�z7s���b��\[绺�*P��P�7*���G�� ,�R~�sN�[5S�7М�:�ln��)��\�0�9����N�u-�n�O�Ksv�����D�qο��
��{���^�뽆��[�q!��f�5%)1	=%��y��D�Wj!��w�X��;���@}V���z�l����7\8`Y}���Ԣ&�JN���(�~�kg*9m�3	[�*��� 	u%m��dɒ�z�J,L�����
����qc�[�j)z�h6AUE3��M�n�����X�s��L�8Y>��o��t��j���Eu;�%'�-��0����P��$���2���m7Lq���ʭ��l�������f��6����㭾�p�v���+~��%���0��y555�q�(�g�:m �� ==};[-@��7�?O�B���҆��Ĝ��(�1[��0��^������a�oS] y�H�u!�;{����$N��*����������\�mo�p�_7:�H[4���g�� ��;)��ٝ��_G`��R�'I�E��F>}vj?�Iu���w�:J*��zA\3P ���PW�OH�.�ѿ˥�N�]\\:?~�X"�d���c�����}�qF\�f�h����4�t�A8�رc�5�Ø�\�0��}էTƧ�z�I�?��F&2"��6H�$�����2Fߐ�kf����η��s�ţ~o�R�i "e����>#-�䟆��JS������v�����;�x��̟粆��n���pY9�t��!�5%��Ep��`f����<,��p��k��<t���'�$1�^ `b=��NB>f$�w����]ZU�|�7����W���/_�n�˃l ���\�j���2,�B�t��*J�r�9?2���i^YQp�<�m]Jõ+���e.�4Q�/>� �--IP|hj���a�Ď�=j���`U)1ᓒ7�
�>�ef��OM%@��_�P�]x�I�K!GA��c�ⅾ�=��.x����N ��1r���6effƟl��Lf�LLC&sm��F�(}r�3*+��(�L�ε}��U a�R9��ӫ���S�	�!�0��q�w3�y��ap��N�]�-���l?X߸g�:��t58�e����99ڥ��9p�W�S@�Y�a5�FO�������7�d���\\����r�P���!�g!����f!ձ��\�S"��~�Hs��y��o[��)���r�j�T�*voh�@���x�8T��ǧ����ʈA��c���!Kh�_*d  ��RW�y�k��1�q�G@6��X>�y,iKb�X�K�}F^�q�������혶$��G�kO����T*8̗Q�@�+h�ސHS-�KJ�:�3:��*L�;�a�,D n���������>Y��<Hv�f�Q�$���-k�?�٢W��R��Ė�u��VKl�O��ȼ�����߱�������o�[4C[-�.3��q	q}%4�֎�J+<x�Fӆ�#�q����a�{��FG�z��V��w]Y�gO��&���d��F*�*�F`*����C� _VWW������y-Z��}��3^�<�,�o�Q<���m��:�<[��?6U�H��F1��(��(g>���M�?�a1�'����;gTV�Fك�k:�u����i*���ഛ�cZ�yLG�/$�����"(���D�h#+����|KX�JkP���Q��§_�f>�/���r�$�w=��Tú<=f&�� ��"�#e���b�2�7���9`�Z��N#8}5�_/�+Q� ��*]��(��R珧���EA� b-s3�Hd5��:K�25ZUHh"�m\n\87�[(��O��@#��'+-#c�2J�*����4��&��h��w;�J�6ۅ[�����8�bE?��^bo?�,V__�B��r`b�H|��
Ѧy
�.�r�v�_��	盔�Ѯ]�gΝK�뵨j��!7�����j�Rn�ٜ�����	�m'b��v�
$��
�*a���~�=�s��?pE`�d�ܝa��)����@�,)_�nB�YW�)����^)j�����Bא;ɽ�k���	T�`�;�cMN�|��d?�������~7���������h^�Gg\��{y_���E�9p`/��_3��H���|�ʕ��beϋ[�[�j6��4�$����i��ܜ땔�< ͌���~����[|�׎����@�;��̞�k��[�"�!I�727;��� �瘸d
�`Д��4S�KYf+5�r	J7~���FR������s�)'��p�KIK_��3M�=/�>�:�G� �9��tT�҅ǵ�VΌp���&��(�;�zo�K����| (V_�:e�e���P����<���=˰H~�;fʛ"ףt}��L$��>j� 榬�T��C>�X�.?C!_����p��=ē� �AP�����]��u��[�=(��^�^����I��U�i0}C{{��Į?ny����r��6p�7ڲEX���G�F�燗�f�Q-`+Uz&V+�A�@��_Ҫ�WǗ�F �&�'�J<�ZΕ����')Za��Q�PtǛ۲z�{o)d�4E(gtJ�v��l��A�����z��Ӡ�'�����A���1����*��7���;�� ��=��\y_O0�f(M)����Ȑh=��ɀ�xd�
�/�mz�RƧgAX�3@���7�o��+����Y50$T��̒[%sss}���z�k�����"$WB�h���C�?�*��L��m���-9�X���5���g�ŋė67�C{ZB�@];w�1�z��&���|3�6�';;{�]| \ �+@�"�<<6H�+ǃ<s�L��De6X�_?vx�c0�crM�e��Hޱ�[$�LfЫ��U1y��q�<�xx��P�?�%�p��{��PZ�M�"�-�@r���"H/�V�?!�N9<�ַ2�hR�лɟ��Ȩ(sc#���e�,,,��hy�Ѧ?���>�6��;p��7o���/ �Q1��Y�4�Q�^vMsB �|�����V���>�2�|9ȟ��Y.�h{O<�D{$�����=c�Љ&�����b�DM]}�,]�u�w�VUqM�qP��m_�E���W�>\�0�݉�E0�w��{�#��?w��f�R�V�t�������{��jOgX��'j�-������E��Ӊ�mFo+*�V�^M�������1^ T�WP��cp��I}�	5�x������V�Nl\�3j���Iڪ�a S������#Y�%WN?ѐ�V��+����xL��xqw�i��Ҷ����̳��W쫢�icp	S.p�BS�Un��R�|+�U������;jN��s��bP��O}ێ����Y2����ADՂ�o��W�}Ǧ�u�x���Y��>}��X�x�u�_/>�'��m��:E�^���ϟ7�.l����l��]���6��R�Yû��m���۳�6ˀ���E���V���eVN<�W�z���j::b�]��O����6��X�~TW{�`�VSw�[����\�/D��(ơ������V���0K(����辩�a0�#?�Z8?zܯ��u�Pj�q9ާpv'�,�P+T�H�;}��sSS4���#('��^�}��2[�H.�*�999���uo�925ȦبbQh��g&i�u���c��t�P�rZ�{ �
QZm�i���ҥK�Rbf�0jB�������I�@!��B���� �,�6y�&���C�ìƥ@b�S������Q�m�m��se�TN˹�[�J^�zS $����)<ɂ��Z��OL�@��"�v��(\���x�W����LQ//�Gr�����G��[}�#u{�����	%���0��+eV�VMC���D�6#mϑ�8t7�3(��5������@Ͼ��т���55���ۣ���uXJ��U@D֩���{��ϗ��e���t+o��yP�}d���A�����s�%^��'����|�ِ�U��sڮO?,��D/�}l�Zi�o��]�%W/�8��H����~�y��g�"��4[�+�|r�-TM%Mc6��R�TCV<�c��o_w��[��(���t�p�hb+�III�_^}���C#�M����Є�Y�K�#��W�� N�~�yh�<М�ڋZ>y���l �A�� �RA"<�]-�|l���D����&9Sw�\�]�`���d�V�P����щJk�n&�Df���Hw~y��}�V���h�A܈,�T��}�b&�Ҷm>]�&iŊ�9�%)��O�A�t|�*��to4���j����L9��b�6{dnL�ʖJX�z�Q�r�(���B�)���c��Z�ص旾�g�A������uuu��ㆆ�%��wns_�xHBO�>�V��P}pTFFFj��t6�h��������T�ng��r�6/|	�2��?��OYUW��t�3{%�f]�3����o;X�y�����#��b
��-��,�i7�w�!�FÇ����ǟ���"�������r�6@?�W(�p�eS�g��_��f��E�l�=ץ����k�Ww>9���y#Vc��q��J?%�U��8�f%(�������) ��w��Ѵ�W][
u�F�uf�2��g�����ɝ�Y�X٪Q��k'�U��Fe���N�-�B�dl�Z砤�饯ǝ}+��]�7;ɣ��Hfh�J��#Ҷ���a ���|�����o߾����~�#}�X�h�o���I�t.���8�Ѵ�+�	�+���rfpwwwօ��yks��v���j]h)Ե^0x	
�;�u�툐�硧�1���SI����PZ>=ޚ�刎��[�����J$H�����LU��T�m��I,	

RRW��b�"q�=zM��j�7z:j�K:�B�]�EG+�Zf����wF��ɕժԈ�zy�������߹{�=|�LJ��蘻U��w��~���K�j�� ĞL���MUe���ٻ�VA��z�*���9`���k�R�D.�ٌU ��Ρn� ATa�~KOOϕ<����%�\�\����*J;�(�6<�bf�۳�<l�k�gt&ill-�=�68͍!ںT�׀[쾾�+y�c�WY�y���Ŧ�91 ��;I�p��u����~k�z;;��vv_^YqI�*D��v渖�8@�	x�A�<�+�ŋ��� �def2� ��|��o\�B_��s��B~9�6�9�U0"���&����R�JKK�����Lq+�M�-��P�rz���i}o'�:�V��޽{�j~��^�[LRPXX���TU0˪5,��3y1r'�f�=j��/6[�����egn�G�</��F(��wM���4<G�3nh����/ETQB��֭[!s��JX�hhhhET�S�/rr�k�WA�;ja�K�r�q�N�ڕN)`���;��N��$��X@����a���S��{LR�\`�[��'��I�|��r�������^P`���A9�`�N�E�*������=��M%� �@Y�ѥ�C#���Oz=�j� �JKJ��	N3M<<��^`��ÿZf��Õ�%p}��$/o�e�b������~��pFL�V��9��V�"2�x�������<��-���7���QG�slD.�}�c���{�G�`�{c.v)��#Z����	� 3A*��yi�I�ni��'��҇Em�2�e��6�5_-N�dUF� �����N�
[jPɉ�2��$��Px�����oh����Λ��Ȍyyd|P��nP�FG���,ژ$�(�����Q{�V����t��V���!��a1+�z7��t~K���m���0rn�u��8��Ij�ށI}D�A�o����D3�i�y.+?���<��PAk�ï���a��bP�?��}*���nT��n���FP�hm��H��ijgoof�ǂ �,/7@��s���5�Y�11�����5��S�+�=)�Aɲ�,�؛6��BևT��CԖ�~8t�|*��*���w��<o	뀂�6����#���ZZF:o��D)ceuݠ��+�V |]Y�r;$$��퀚���DChe�B�y>�/D�y�����R�4�`�l===�es���S�@�e)"����C�j�&xWy��9�045`k�0(s<YS4�8 D5�ė�.Ng'��{	�.%%��*<��:����+��&ZU!\2d���h�����AZ��WI�1�;�v�f�o��Z�V˯6 �hyO(�zw��:@��a��/��@�q��v+2�[ �CjWv|���iӦO3��Q���1�?8J������:��*Z^t��^D8q��!dɛ7o��w�xf�ޚ���ؘ��j��5Ǫ�!��J����Sn��,_̢�ի�����ѦI 6��e8�}oo�N�Ү-a��t���_��ca�8���	�晱�a������4�}���!A����<��U�Ǳ]]]���y��w��Cy�RqE`����l���36Tg7f����E��l
���&���:  ��ɒ?��2�&�8��!����&۶�d���ا�GS�1��9�L����e��x�H@�u]h����G�N�8�D%��#����.9�v�e>mG|B�Y7<_{Bt��ߒ0�*u����Qq��á��pA�𖰣d��H�C@Q`,Pt���N��h�S�=YN��-$x�V�;��EUf�ΔWuIGb� S�j�F��4��ܒ��]�� ��(U � R�hU͟C[���S��!L��b� ��q��������j4 �N6���7��xt��pE�ޓ���a���C2���J�����n7�<�U���9Z_1�c�����	�PD˜<�-Wn`��g�wP"�8k���O>�jW�h��8��K$�ԏ�߁��sMT��o"���	�$�M���f<�|�\nL�ɱ�b$jNЁ�ˡ�t�9a�ǞT�m�H��i$k~�H�g.��"�4���17n���I6����o>)>�l��͕}��|����x� �ٸ����ɓ1MMM$)��n��|6�t��Q4�D�TA0/�r�'��.Į���_���Cfl�����Ty�A�W~��������0A
P���)�."������"�Vq��h�5����#�\!�����u|Yҏ���j�Wz�]Q�>�8O� �ךʫz�+rk��7���P�t��B^r/#;;{��`�L���S؅��Q��Թ��jXWU�j��{��r����k7�ő8ן��"���&�9��f��N�ɵ�-�[��o��ͨ�NUUH��!1`&�<
c�W�M�$�w���m	nBJ��|}���D��}��7�&�R�b�>DE{zP�/�h:��!����_�Z��"�0��j��7P����c�ջ�ě&j�~�8U�_�;��~�yPґ��J"*�����h^Ӻ�0��@ظCU�HK�s�旹I�I�����>Lz/��F ���X����2(��:	�����@��߼)N4O�Eo�ݸ5��@~d���Y 	�f���w�׶-���G��c �������vm@1{��y���������ܳ+��؇��Xo}���D礏O>�k���ݷ��sM�2_!��T��i���<By낳M:��ও����0�z��Ɔ��`5j�#��
Q��	��m�^�M:@���(�@����h��g�\���K7�) �/�k7߀L���Y�*"��7�rOw/���Q�����=z�TyB����1�oX��L�UW����A##Z�f��9�����G=|�EO��Ɩ��vS���sՄ�g%pi[4�/���G�7w�e�CK�<�ӯD�Gg8
(��*nZ@X{�ӧk�}��\��-��򭪲��s+�ړS*p��J�34�KE��w: a��F�?�a S;~;o��ic?��_<�u0���Eԯ���P?(͛9#,���x�n�V����or|�EDE�5�ֆ�䖏��F	h_R ��C`XYɧϵk�Y�$M��t@/����Zû~�����{m�[,�!��m�UT|heM_VE{qBu�^'h���@{�ln�)-'�-�K!��5=t��ܯ�7;���^VV��rA%tl�U���>E8�<�H܈J�e��r?:�
[C͓(\�/����pՑh�E�cǎ�ŝ�a I?����T�{{�������'x7�����i��"���s�~ϰ����}R0�c Gl�W��a!������tt�[���&�߯�ߺk�44"��)(�����ܝ2!�T�}#��,D��${ X={VZ�7��x�&k�Sc����L}�=y���,��:=��O����_�"�����G"Ztb��\�m�>�>��v��	������!�{řv�mio�!ع���l��n��!��^^������ؽ�1�TT�'G:ϟ;W�ݲ�)�^���~����2�� {���er�~�����a���;O�f�� 1�n��m}���\A[}�^���jD�b5�0�¹h��{AmiF+=f6�21�~���)�����5BY������2ؒ�1$.�#����,����_�:I�^���YR�I{���B"����̽GE�6�~�0o�=8ߐnot^����]n��"H�*V�;\��b�|��)�H��9�"�'z�x�v|������/'��_ru�[������8���F�̇b���S��T(&�K����?��R�r�A�n�H�Y}�/�(�$a��9���4��������[�|D?{�C���q	=���	�{��Hܒ��β,���| G꣥���_*�B�7��⡣�<*��,"hh��ꚱ�Y��@�pf;�ZW�������U�! �%���0�/^Ƥ?4�!c*fz�w���ߎ@�������}
R(�V�j�`Ծ B�	������T8=>�[A���sZ��h��t�^��s�=�D�QȮS��%�T~��t�����lvh ����N9��1n�u������Ӹh}��-3�g:��FۍU��M�.hK�(����KfA��k6m���{�TR�6�up5�����ƢFr�(�(�]'�h��pj�m����h�����bB[,�c�
�9}l�y�_��C��و~� �RA]Ą���ui���?{F�q�tM����;��Ũ+ܶ rm� ����� ��� l��W6SUy�b�\���DZ�Ԑ6p(��d���~N:��0�Ҁ޲!�@f�|�+R�=���A9nbf�긨�T;�,�l����h�
-��"�� �7����K�eP��RQ�8�O�8���%�P)o/�� ��fYk��L݉�*v�`� �����I*��"T	f.s��q^�c9rǒ���+555�ܜn��n��^�z�*Uy7f7?�Rq�J���!m�%PIn�R��U���J��-���Z�I:�]%���ׇ�Z�^���J-��B�,���vK��:դ��Br�X��Y| G��$��&�V�K���
qM.p�]�T�U�����4;���aґv�C�-0X�摦J�!��\�h�D(�F������:Z�0���9w觽x��&r��~��W[�b�o����2�u﬽��t��4���7H3���ٯ����廰��UUؖPƏ���"eCD�*��v���r����e����2x}�/h��.�Cc�aqޕ�GRԚ�8L���s	�dϐ�� ��V�2��IJE][t+����qe%���f���Gϟ??�R�Ә�赳��8z���(�������㼯��@p�S;p;!�^ǬuF�&��˗r�XD�
ѫ W�����]{͑�?ω!<.�*_���I3��͛��O8�"�D����Wo�fgd�}xK�ѿ��F��R�Є�bF9�Gf�NMѪ{Ƕ �u+)>����`�˃kײ賴O��M��A5��1t�
,����!"J���ns�9��ȱk!D?s&)<2�ulBh���+�G�H>k����[3��X���f&G28k��,�e�.���5�7]�te%�$�ț�^�ƾ� /��l����f��u J��1�@!���Rc3Z��X�/�k������h�n(��]%����}��>М+9>�| ���n�FFF��p�W���k��q-�5�����YSW�ìA�b�@��~�Q-777��b�L���\�Rm����&���Bs6*v������9yF,T�P'Uq����O���yN:8��NKk�g�
��lW�G���՘5��E򷬣,������ds[�������0����1��o��u�H�߽��_���̌H�}��{	^/�ι�np��nh�|�������O�P�cA]袣0b�׈م��
V���4�\�~����X�R�P��<��Im��>�N�"���^C�~hh��3��d��W��:�}�x�kjD]��l�;9w����.��@��?c�回�6�Β���Z=������ΤAȠ��TwBu��Y�.���4���q�Gi{� Ru~���H�I��������伯�ܼ�ҝG5�T>�놠�+?�R�]���艶h�$� �G�j�D���40Te_�3&}�o�N%�_!>�Wg��F{���br����K6���}��ᶗ�԰P��U�B��~(��5����'6±�7����!�AE�^e���t�*�j��K@hؿ����F�cd�4��Pd9	|�
a��x}�ا�*� �1��TBOeU���6oMj�O  }��e�S%A4pd�Q�΁t�ݮ�ڥ�EpC�ѿ��ű�5���?{$~s`5�ǐ��c�v�8��:�R�����jjR�{e�n�47��S|��%%y�����^5j���܎F��p����S*Z���[���;��zC��v����*�Le�c�u��iiκ���S�~����wTF�
>=�����D�}O�O����m^\�v���0�3wwE
�����P�Uh��܇׳ڐ���־Ҕn�V�3x��ܷ��g��c��C��4UN?�s���]G.�?��_6��n��`�B�}O 9��qR��V�dR}/*E'Ɛ�J�J�4�����	��<�_�'�f�G~��G�����O�F�m�F �j�Z�&�m
@(X7A�Ъ�l��J���egO��`&�ܜO��!�z�B�ugU4"��h�TV,i��QL2����Ǥ]�}}}jّ�
-�䢢$�=s�cI��%����J�sݛU����J}>v�)��pA�1�y]���I�rJ3=}���=�J6�t��ܓ����3����'�!�%`lz�����D����a���!@���ґ���&��0A��Bp�ÎSo?�f�))��F�� C��{A"0�u�E���P��/��	�Ѵ��׀�| d�|�[�Q񻼊v\j|�Ύ�s��!	��ϲ�P)�N�c0�5K�`�HDP�����|(��s�9c���WN��y%���J�$�����"�*/AD|M�j�w�7j������ݞ����b�L�l6"���:�	�%#Z�����(�0�U�F���0����~]�믐�cц6�^�4 8��J�Y	�b ٝ��F���e��&��X��4	��sKJ�p[/��,�K�v�p��C{�^��� ѽ�G;&cI��ٞ�`Cc㻸x?ת�mnh��BIՄU�J��r�B݌���L�^:A ���c�|�}�x�f��S�����;p_�S������|�q����+��+z{{�~��Zm��R�~�:���˴�C�8�Iq��T��<6��'�_B&�4ѻ #c�i]��0��ћ�g�R�A�R(�X��yK㊐���ʢ@T%Q#������TG��,�M`������F��K������L}� ��bFf�Dϩ��|�ѿ�鞆FN�9�R�H�$�`K>��?Fی@l��#�9d�ƿ�7���=G���Ǐ���������{�5�c@�<��gɂ�htt�$O����<fiIbef7�+��=�i��'ܸ��F x' ��F��ы��_�� �βqla��Z������g5\	�8S���*�;�C��ܹs@{�Z����/ßf�O<�!������@�zL�ihBj,������z���&{�%���|�L�R¾צ�	~� �T�
Ϩ����od�K8w �vA�TY�4k��E��!p[��s'.dc�4�,(�Κ���|VA��/��+;-[�hA+���z�hÓ]����m"��fblg]�D�^� w}�����0��;}a�z��ϳ��qwڑҳ�����!jN�3�PE_��=��k�gG#�b�-���z�kc��WY
_u�����AAA�"5���P��\j-Z\��ڀrЙ��C��/ӆ��m�W~���v�+���b�jh�O�hK�r�Y����V��R	b%_�j>��F��ޔ�~��y�.�<���������Fp�n�h3"w�=���4#bu�U������N4O*D;5�{��x��̓J�����?��}��l��l�*l�
�zH�	�� ��k�r����d|��1�^�tx��%K|�A^u�B�������m>�	���&��
��]�̻�Zlm*������}�ݝ������Ƣ�SR��@kL���%X�M'���/�	2��J_��`��-Մl�ŶV�<n��,�FЂ�S����6��J�W�0"���'~�BnBKW�ᯁ�~����⤻����N��~�X(��w�A�H��@��ƶ@�啖������$��b�T�`ccc(z��5rD9-/�2%99���E�sá<4�]a�h\��m��S�hΒ�lE퀐�����yF�' ��Y����t�N3�9�'""�r�Kx⡄�goo)�~��>f���<KIYq���1��d��c���������+W�`/�'%�]�@\8�y�1���AMӱd� n�قj\��L�� ���YH�����T��7M�362��CVvG]̶��k7��"�(i��~a-=������x��OO�[��0�? ��V�\��MY��C�b����$D��p��8��卙]@���{���t}�{�x��g��B,
�8/��rBv��G��'ћ�t���� �(ĳ���_y#^Keu��qSX�9��;�c��*�h1
e�r�X���#���)�!�j����df�l56~����c?���?��#j���H'���ߤ��P}J�B���Y�VP.v�v��,�1��|t&lEG�ӡY��w!z�Y_�V��;T��i�o���BuXS����ڏ���Q�`�H�=%5U2,�Qo��Bk;򗍛	D'�@�N%����vq�Xj��nVR[{�Gj�a2���(�������ǡ�N����7fـK�߿ע��-5E4ƙ�*�Vnz�Po���x=�3����,�첲2x�-.����eo�R@����2
�+Κ�)����bxr�K:N���ڕ�� �����������mS�{�ҕ�d����Ay,������O�Fu�eg�-��Eo!��\QQ!��e�W�Pg�q�����;-a//��o+Z���xN&7�>�}X ���S̲ɰ����h<ݾ!#�̘�VԈ_��t�{�N����GR�JC}g:0�#.���UmoAס���9�����C�H+)n]����w���&�;v�y���v�G gd��3�ց/��l�������z�n�T�P%��`�'M-�C��@�r�[u���3�Bښ������L�����%�#��cA ����M��\��qIQ)K�JHʾ��5%elQY&k�d�:�V�5{�qJH��K���S�X��${�����t����>ק��4��������y�!��R�m�	�~h��:|���A�rj�S�T^7.����˫M�-���a� �O�2K�"v����7F�t~�D�	^�P}?x�16��!��My�_��,���{(%�!Uy]s����#�������4z��`z��	t|�l�c[1����w�L�u����Q~Փ�"�.`��a�aA�0m�;EZ�^Ye�^2�hy�S`�2��}n;���X��1�����������{@��q@��ՌZ��B�i�J�W�3���yf[�>e�]S{���ֲ�[�ڨHr��In�{><lq��L�e���}<q����,���\A�E�_\!���Ӆ���;�t|��@t�I���_!Q-XC����o�ޤj���^�-
e2����Ѯ�3��$�c˳��͛(�d�e�=��p���iYY���R�;v@͍�d��O�ty��k=�ȶ��>�a��	�cJJ�kݕ�	��O|Eb�������g$��)�W�
c���!�� �Z�x1����א��'9*�;��wB��*� ���	;�s���I5�y���u�6/�m����M�峗��Ⱥ�5�r'555|���e�R��?�Y�^^F&&&Z��NbO��2�V*A����03��e���|��v�LB{�.��j7ev�  �_P��e�9,a���vv��i�t�g�t�������2�&e[�-�pq�������ϟxh��~K�ī"_�8v�������%ܴv�q�}���RS?��|���V����!(�pA]��9�/J@�aԡ����B�'���H
p7������H���P~�KK�TX�lon���?�	��ڋ�����gDq ���m���w~�(�����`]�jWր�nq��^�C�,���T�]�ꏱpǉp�	�.���sߜf���p�Z�]�b7�A$Wj2,rt ��Asm�گ?�]Y�ɇ�����[�tx[����}�P��x����"Cu�
[l��E6�ɌUo��=��,)5�:���
�F$ ���:����Õ#��?s������Q�3ä~�'Z�o�%a�w����^�D��;�-��H6��1)�Z��nD�l�;wP����=<�>�~�W9=�r�I&�����iA��P[p��g]����	��i��3�R�p��E��>ii���Smh��A
~��8����J��SN����}�/¡���5:3sV���и_u��­9��bI��3���+�8���Z9�E��fX)�����;����եw��?����Q���v�}�k�.p��U��)�t{������m>��?�6.�E�'Ϋ1D�y$���2��w�#MM_|��M���!��#OY}�$q��b+���A�"�M膖���e���t~�6�&4��M4�g��U����jx�θ(u�Ν���P\K�ƹb�����h�"��<9[� 8˵�C**�yyyOJ�GG�=�_��5�`��t��<VY��u>��ǌ�v��\oooQ}�<�����<fnm=�1<VYX8˥���xSw�[�n�B �E��=/UT[ۡ���L��������ϒqA�\��@Kծ�]�7�m��Pɡ���Іk���mmzzz��m'�R���-藣��̰�%��߶� �l,��^��G�
���"�%���F�����KݓySQ�˥A^_��yS-ls�@��EQ$
�%@�F��.h����[h�G-E]5�X�uS�m�Q�`�S�1cQ7�;ޯZ�n:r�*;�yG3D���	h�}]ޔc,�1 P��K�ɐ��b����3�<��[m������Q�����.Ղ�/���M78�����ߢ�1�$EG��z�@�@>�f��Ǆ����Nn���X��MCGggۗ/O�9i�Yo��C:����11�(䡽H�E
tq�LL璲˷Q���U_�}�xۇ��m�.0B�����T'�w�0�6�Җ�s����G�kfv�&%m�Li�>w��h�S�����CX�7�!�q���,�O�?rn��I���mm�2qC"��r�/��a�,��ꁯ��5��&31� go�Um<�l�dõ�k�]�r�g�$�d��l���`w�EBh���@��t�u�Gߡ��+Eee��R�u&|��O�5�C�O'���f|AoBd���	ཚ�W+e �j
��ΫNsUT�����3;,g�J�\
������EQ�*hb�cUr�Y%9���}���t�AX����E����׌q����`�|6���+[ގ�_��!�
3]=�I���,��Ȁb��q��Vp;�����J�]f��b�>�AV��|��e�FK�����*�3�C��ki��b��}��qk<詚T����Z������}���`��T$CX�y��b!'/��}��۷3Pڣ+�^���bQט�mѻJ�y6��I�>'''2\#ഭ@�\E���m1�Z�~�j�)��a�8��鐽��'�?ߝ�:=�f X*Z�$Q� 
��:�"e�o��Wm0�R��U�Ob<���~/�@�pCu]� ��#١�+�
f�#�E��D8ޔ����
���@�Q�?**//��xs���V��e+���5i�y�5۷o�����׾}{]jz:�n�ά����Ύ�#fU��:YZO�zj!�`���Ǐgj�ӏ����[TW'��%
Ԫ��ؤ�.��MP�y0j&���R�d2�^ۦ�ΐ�T��	z��E��p�ތlId������p�(�v<&&F�):갾CP�E�r��K״�[�cd�.,�U���� �v�[�N1qS@�<�ua�����+{���g�ѧ���/f%J�2��m�g�%��"D��LLM��d��Ǻ�@���t��>�ˊ��X?��c�@9�"��S,s���|�M�@l�舆K�Ū���� 3��_B�����.���>hd�w���������:w��������i�9t(j+*̅��&{�|�<M.�o��z�e��A�p����;�6��b���V[���dFu�\�̭�,&�jp����S�H���Y 'p�f��o�P�˗�8ݱ��D�P���NL��kuva�P��D"�����e/���D�����N?`�B�i��$�F����8ArQuu����g��9�R�6mz�5�KT'^�3(H����b��;�Ah����>��Jc����t�(����9�qu�ӧO�ǡ�m�0�A���i�%���R� %�/���*��uw'��$g'(܀ܣ�
�M��m����6�$����x�!D��������q����	\ �͛[��a��vӉoA�f]�&�ŀ��,�R(�ѹi�U�u$i�c��OB���Ԉο�~'�rN3����Rca����e0����h��!����Q�ﺈ_C'�=i���>K���w���Έ�K�����L|�����}%K��뎎��?%~�Ӊ�韯=����ǿ��Kv��+���:�op0y&��b:��Z홐�8�K���e^7?��ć�"6?��ުz`��������@��Ʈ"ss�8�F�Ul-s[�*�!���Xyzn�c��09v�)r�U//[�h��C������pH�fT���"�+x�4��C/0�p\�+�nFo^�����^����=�7箩<N|��nu'��)l�V�%�����;QUTZ���	�E:�v�ny� Hft��))�\ܔ7�}�;�W�'�_>�%�<d��ȼn	u��ϟ>_��	~�����Ç�WJ�6g�W����lP�s
��K�켪!�j{�S���Θ�0�h�ߥ�!�S�P_���H�m���3���6u��`M�1�4��[����������a�o+�����s�L����P˲ �ݨsK�v}I���pŜ>�6��c��������n�d�~���w�-CfZ��;���a���������5.-I:Ar�$:jnnT�_6E��4���Ҳ��9�o�:P^��,{���򃈽���7~T�9?/F9;|��^���^�ADz�{�IX�F��6 Xݨ [N<QQQAV�)�����8%� �0 �*U�^>�θ~�r/�n��O�-d����p����btQ����mހ�@�B*	��m�����)c\�w�b"�����TH=XiM{e�t"�x̂n�������� +#��[u�����5�Vch������b�Z��zmDJ =1��e����Ր	�!�"z��@,�<Y�ZFb1��ja�?R�:_Qv��AV�>4�
�'�@�dj�G�b6w�/�2�<��D�UW��׎�i���ީ*<L4>��(�����o5��uT����p����Բ�[_K�$D򖭄�U���<i(��-Snn������l�~�1��J���f��a���o�����)h����P����ȿA�����ā���\�&���ג0C�.(,ܾ�R7�gb=B"\�(�5��=���+��k�6	�-���S?������&sD��_��<)=��*�`�C ���KBo�_�AA�?��*����N����#�u!��S������[��T�L�'񤣏K;�(�߲����C��M�	��-�}�� 8���}�W.H%E��V�v1�"�:��;����W���B��B���O�CU�u�R��
�k�'ؙ({�lw��h�1�Bᶧ�/�Tx_��z���*������7\<���XA�1z�?������dDe��~2B(�{�A�"�
}h��B������E;����~;|���l��!U%%��މS5uլD�w^�fU��j�_/�Y���)�D>�YUC�X s[ ���CQIvySV��
C�z)n:��"tp`����4/Ar�玿w:Rғ���������c�X��Zk��@U��gq�@���{hf��,��E2PΠET�ٲe�ȷo->=-�i��lM��H�F��N�����^���
�.��.�%�~��g~�R�ˍ'����ޓ3nt�t�*��;F���Is�;���W_��A���0ILcZ��AAveh� ju�O��D؋/Z޾��)�}�p�B`��)#i��l7j�LN�\��:A��Z�s�<ٜ�b*<:�d+�V���S�}%���04��H���v}X�s���pV��hL=�� p�3|��� �`$Lʩ������Th�l@D���b:��th�P�'��JN�6c)tS1��^!�ϫ��/ΗO�.����"3s���g�!uV�C���h)���USCƸ�UUФ��c ��K0rX	���o��:S�{(�h�j�g��DFF���u�۽�*�����g��|��Cvn��WV�����g�rc�!���1#\����r|�89�d��˭�y���E���h�
�=b~�WNEf�ޟQ5$� sB�Fn�Ǧg=-mEzh
��E�4C�� �C��I2����*���2���$�yۼ*o��PYع���\��> �����W��D�� ���qC�12��Vr1�����Z�t �;�P �R�Ml���@2�EN!4��~�m6+�-v)�t�G9��3�Hwv1�ؒ�L��2���;��n��!C)�$����7aa��K\�I�S x*'�.mIv���g�c�w��8Q7�0��,�D7�B����������~�"�g�6b���	�@�� Y�td�3e��d��d����5�r]H����f��O���7�\<���y�Һ��I��E`�R��w��E��̦)R`]�l
���в�XK�19���t�.ߩ��$1�D1�p[�SF��I�.�f&X�Oh�'��BF������>�[��C��$�p��|��	fɿ�{zzV���(�]�6D����I�3�r�{I壣�6�ɦ2B��N�-�_�t��+���y�5�Jǥ6��\��H%,9�ə������~ͯ���;]�6�X�^���Ѣq>��e˫��]�M�茞؃ѫ�P
�P�� �j���$� ��Yyk��w�\m�zt8�I�4#�8��.���\�N����I`²�2��>�%k7D]*� ��G+�PK���^��!�pN&S�+��.�'{�_�jlU��L}:3��`�4��ji���1�ӿL*n���)��.f��6(S�G҂����qbFVb|V־��������}Y���U���:�7���-�u1�l�����Z� ӪU�K���}��;1���G0�g�4�,g8���J�g�w�/��o��x�~9&h<MU����G2�YC�.�0�c/ЩW�����!W�f�d4�����cV6ciiia��D��G�8�q�_���䝜��K�F���[� �<�~���+Ҹ͇�dEDK�D��&wM������$E�e0C%H*���_6��^~qg���a��ɛ7o����g�R7���O���Np��1=��f2+�����װ4�3��� NPH 4~�����r ��^��sLC#������k�Hl��w��w�^�j�Ї���a���T�Z�����Q&�n���(��Jd!�cG���.v�A6�ə��j��.��;@K������z��v��ϴ�3��$�j��נ��z�(آ�"Ѳ���u��v|�u7qX�����z�C9݀��T�C��l������ûS�8w�2kim�G9�Q�?,8���Ը۷׹��4���~����:n{�Ϣ�G�jQ<f�����P�`a/�LBC�\�Z೛D�їM�۝�C#b�)̯,����L2Vn�B��WL�� 	���c�����\�_��}j ���l/��[]Y�8�5<s��&�2)�L&b�
����{���~�j���Ӥ߿��y1�o��,��P����71 ��'"[�r(�?/'�r(-uؽ{wnccc(���ʌ����{���{ƼWǰ� S�F��7�ZzY�P��������2t��」fC��"���N��n�l���]����ig��Fՙt��m]{�c�L���n������#k�N�鋯Y+��j�V"��8����:�$�F���w�Kz�%��;̆Xwvv*u,o�a�\)}����un��,�AyÒ	r�:E�gT��zG�*�w��w�d���T�v�؍������&y�P|~���Z�n�?kP`U0�%��1MRlm���^>#��u�����:T���Q��[f�+�r)�I����@�/�H�j�i=>�2���Y�F=�e���g/f��0;���L�8gcK٤9O.0K�O�?���W��4��������5�O��+*z=�� ;�:��������![,C�	J�Z��a��U�h cn���b4��@5@ä9U�۶?�k���Z���`�+��5O�jTx�L��^�;�w1�}�=N���t595��;�oJ��ttj�-�k��9�[�i�����w!.L��s�Z�v�~��Xj�ܠ���%��s)>�T,T����R%��I���4�Β�zex�K����R
E*B�)_����XC:�A�׈d�7#�e�۷�y|Y�,���ˌ�Dh.�n7SSK��܄�MM��=�٦�e��p�1�BDӥs����~.�	���$=̓���gD�ӵ�*[����^e�xN���]n��B�6��en�ii	�3F�����������JTgo`xY��;"Ld����-,-S;w�Z�FJ��������~~�.���T{u������1εp2�3)��2����3�l�'��e}��뎨��WCy@�-��w#w��.+^F^>��!PVY����eo��0wH�G���u����s��r�"�
�.//�È��~1�$z�μ�>��s��1�<���i���M^EnAU��D<�?��eww��
�h��z_�8�##'��2>��%F-������fl�UÜc�l�̗�f��2�KAsV��I��ܓ<w��6sKK���44}1Z;������322�[�[�tA�]��^�f�iF.W�5�:V��w3:;L.*.ދm _�x���= �\�*7����O4��N�� ɝ���Y��q���][�� #�<������K���σ�ysG�s[V��r�?�q6�ĸq��H�<���_��N��-7��)jY��>׫��= `b����� z@}y�� ����m�f{��Rpx�T�E{��P�MR�U%�#�F0�L��/)�sHEC���\Y�V�I�Nk�t�L��d�i�Y�kgM����~:��B
��)��8��ɛ���PH%��;��SߜS�ֿ����	��	5?�S,p�$7�8nѻ���	I�h�F�Of����1)t��kҰ��N�9���k�T���<��K2�n��h*ıu�ge�޻��v*~[s!��Ȼ��E���:�:ׄ��G�!��H_�rAlll�AL����j͓�e��(Š�A�c����EO�m\����4��)�uܸ�g�;��>Hs�*#f;_��N'ϜKv���3��/�x|M��p�ܗ�M��
�k�����ѤĔ��������Wp΁h6�R��ك\_	Dd��q���W���j�R�i��0��"
�l5��|q8��{n�����}��͓G�����䍻'��ů���u��y���������CZ���(}QJ�R�V�O���9�����ﳐ���Ѵ	C��.��Oh�v%(p��"Hq�
����zV��$VV�5�CA�v�,$�7���:�����Ѵ�ꁣ������,?+�'��P�r�����WY���@���/�Fv��27�L���j��v�c;3R�Iz@��|==��c��а㪟���ˏ����8���¿E2����܄�q{�X����a��΢߿~��X0�`O�)H�K��~�ɝX,#�h?�V����L�mN@���p؁=����v�v�T�4c�����!2�,���X��+c�[�Pn��G���|?�Z/��t����8:9��tP޴��h��
z�6g����'(E/&@��b(sh ��FmY��mMn=��#ﮔ���pɿ�k-s�2�0�{5 �2D�=٣K����	��M���Y�Td�̖\�a�hr��=ep�ر�G���~LM����{�����l�`� �y����	"r�N|?�Y�8��c��/#�$W*�_�m�;=��S���$�ʹ?��ў@��k����P|r$�$���KHEI��<.!�o�W�ou4(��\"��U�/
��WR V;88ܦ�)cL-;F�F�n��^4/���(f���X6���������4\�rhF�$��@��n:�o|�`��+�Ru�ik�㍟f��G6�"�fbz�k*�����i�B�Ą��hHk���^Eee�J��(hh�����x���Ȼ��f�[u��B�����>he��{�wl�ؚ�'�Yņ���^0 �Bj�)��m���Q�2//#4r�a�ӕ즫N#���!~���M��˿�KP2�<�B��Jݣ�t�K�� �����f[S~߮d��� v�X��K�y�#�=��}��D��{���"��/��M*)�J��v	���Ivv'(�",�7lk^�_�N��J&�>�Z��$��_Q�bA�I�W�l�W��x������U����u��u�&W����.Ɖ_�Q9v��0�ˡ�O4CZ���X�߶��\�ꁗ�.�"�)��yɅ��us(�o�fԝϻ��k�cUS�
z��1�f�$5�==/uo����	����v�}|<+�ͪ9R�O���[Y[�k��f됈�N ��VV�?<�p
����27��'7&��.�����δM�z=9l&�(��x�c��'����Z�Nn����0i���ׯ�$�#s1��o2�{�MG��0�P��S�G�����|l+ҋ���E�8 2�ӟ̑��5�u�32K� �]
�mHI�źs}r�W�0T�ռ�I�C׼&�qh�8;[�cz:���t�l�^n\�67[����oh�d��"�!N��@���_]8���&�����T$*��a�BX�8V���,��B��Y�X;������Z�6�5n�m����E/���pwW�	��$�m��{mw04y����K$6^����M[����w��fB��P�,��q�4'Ԥi�U�Do�>p��v���P��~273��Sxߡ��ο��+P�9����!uUh��!`6D���?��~Y�q�h�F*Q��Ka���ɐ\e�ph??�h���}�8�y�8@�da��G
����0�}Q�3�S'T%����D��ʢ~�|b!PG3�#�?/i�B�@���h�fy�%j����
$˴?��h[�ǩ��FT#ğ>KnG%����-��X��S$Y�^���+Ի��P�L4�=@6G3��� FP��2{X�U}hǿ�����)�3�j˟�"݅�h7���ssGA���<�*�OQ҉W���^�STX��9E����T'����<��ğ�0i���6j����������9�'S��QZ>/��� �9p��)�	D��!�ݜS#ny�W�u��0�fI �5{	�����<�wt`]M$ذ��lܡ��A�� H��a�����c1��P����_��d"��ı֟?Kn�J -����^ԍ�"j����	�ի�U�#�q��1C�>T��o�����SiQ��G}s��x� $q�RX,cw �1�mL��������3k�����#{�AԎ%G+Ŭ6�ѭ�Q���+��1l�"����m��(gS���Ő��l�ǎ��N=2�}����^~�'uN�@�رT@�	�h1��Qh�tmva�Y-��=whz{����L�(6j��i��q舽Um��2{���Lc���t�.F}j����؏��
P#s!�_�B�|�F��_�:R��r:,���[�Ti������i�dkk�	q�tү��J�N`j�8'j��SF��^�S튜�S��c�@���p	3D�"�h�R�m� �5'±����v	��2��W�`ћ���H�Ygg����h��$/y����z��R�[��;�@4\�������4^�yq�;�Q�Բt�K�2q��ܛ��]�v��]�t!?:�p���-��y)��U��M`}��i�%K�����ݵ��1%�����u����h�>al��cć&cz}�f�p�I	��:�W/���������e;���c�D��l��JC���Qޭ=)p�n��9�>-�yT;�/�2�R6)nķ,�ŧx���Z�_3��RF|ts��������z�i��`issū�Z�(t(%b���^UYƒ�2����wg�
Qw*T�v���[ڳ�<y�dr�WuC
�m�-	��� �Ӛ�R7�
�2feeV�v̰:�I�T'76����B3T�g���\��c�������-y$Î�yh�XX[�Ƌ��2KB�i*t���p0O�*�.��%͝u�~q_bo�u������q�CC�d������u[�.s���1A��o+�`����xm��`IEE�l�L�c�$�J����W����O�x&�b�����?M�N�׉�*�J���3��G��e������k��Y�LF�D��̦D�>��]���%=�Iae��[1�*�<������@�ȥ�!Z������� x ؾ>��E{�Ņ��8I��:>=Nqx���`�)�q=xvM�e�e2y��>O��L������?�*�j+�E���Uy]Cпx�d�e:zkH4�yì ��nqY�C��R$
���^�݁I9��6mB��N��u�B9���&]�3뼔q,^��ʹ.�"�yX)f�jo�s����q�&y������?+����xF�*�@�(��
�f�̬��ē�Ca]��?����CS+�S�AN�N��~)�#f8�|�'lq7�\Df���e����Ɩ"ֲWJEz�Z��Q�`3l����#����ₜ܇&�U(��B���<��D$���_ȩ�����fY_�r�B����P7
� D�
%�}����h���Qh��OFȯo������LLLF>��|Q���P�y�qvѯ�-�:g�2���;TQ���U�3K��)���XV�.[o�T���U���w�6Z���5ۿ�m���b��`ͯ��G�Ï�f����#�Fխ�W�	�}x]�$(k�dDgg:�����`3k�V�WA�=��_5��;8��/��A���`��кF���s��X�y9��x�M�ё��-A�5��ZA��
-J�ȵx=�oK4V��R����^+�}�e�i��hz�����މ�j;nO]�xq8z*"\�_a!��AN{��Ƹ��Q|o{�����`q;����%7	x�܋�tz��!1IX�6�f�}���$S�8@N���=��i�S��V.��Pq_���:H�۷���O@:%--msjr߂Eq�8~TQ����4d����Gp��C����x��S��j�<jҩ�C9Z� ������/�����o~�q�� m�O�4E���Єk9T��/�[�~�s��?f�T��r��W�{��&]l�@{&q0o����2�u���Aǫ~��q���w�'���VWW#�@��Z4k�۱��A�-�F>��0�
 (����_���q�Lڗ���Ek������+���E�F��GWC�d��"�xrD����4�����ѻ�E`i�̊c1�U5�J�xJqF�E�1������g>�(�'�^]���_�.�yR��bc��MOT�YL�,�(�S���/��]�P?���m�h����k���
�����v�9�2ơ���������
�z+Kѻ����8���>�i���yr����2?KB��v_q��մ� ��I��i��YvM00ff�A�ir�����3��z4���5���lİQ� (���*�Fjݼ�6f����4>�T|�=ʥ=�ekd�J3x�U��hc��mf��']dS��!��4,���ۮ
���z�N�y\���yU祜O���h?�W����i�h�eX\��8���zl�+�:b�ò��fQ���� �WVJ.��0�\�jolE���Xl�js�R�ǂ��+>�Si��1�bu�k!'��߾M�=�d9���G���MvF�ˢ>�R^N�
��Ц��jҾ����qwr��}�(	�Cǖ?^�eH\Qln�T���x�&���ݽmv���0�S�+=���v����v?�Х�I�#c շGX�/5X��5��iXXE�0���@�v 2vii�N@1?K����(4���x��K�o
?�����KQ��zҤR����2�|�ӆO���Щn�O����J�����.���ؚ.j��P���}B�>_��X���g��?�qddd|�(�Vu��:��8�dT=����m\\��,,>��[z��[��v�MSd9��\,y_�ް �S���1h��g�Zs�8�˱M����6pT�=�;H���V {��O�"�ɿD ��yu�6����?���]$�����B�r�:͗;e��z��b$PS�5����w{hu%��6��i��X�k���<�X���U�(�q_D�/U���8I@�Ᏽ�r�޵�����紹�{�M���J�E�����:��Xj{}ɚ�c��GS��χO�=�=闞�����k"��?��@H��T��Y���q�mW�T����y�U
-���Qnl��l�ws#�
p���.v�tJ�c��!���IF���۟$�y6����M�L\�|��Ea�9�k� l3���f?
i�������Q���y*�R���7����R暵Y���� �i4u�կ3s�fɿ�|̴�ᩰ��:��ֱ��k�lͤ�ß�� #�k�V�=+1�0��q]��~V�r*j߉��7���ky3�ZZT�$%%�HNHs�=Z�'� K���'��)��z{��с�D�w�=��R�!z�����Fv��+�W��ʐ�:�e�ն�vJJ���x\�k�u"��'p���+\�+����(�aԳ����+�T��F���b���0z�Ə8��"V:
���n��C���l'�5,����	})
J��̖G[�6#vs��3�%8b������v��!$�2M7�˼����X�2t�ʾ�&�ڸ&-�!�k>���wa��
�(b�
V���6
K�.n!�<p�Nz�3	���i~�{�́}J<4�6d�ӑ�V{�P�_�<5�J`-�=��5�ɜ�_�<ئ�.��|���m�x�W��DB���99�X�&Y/O�!���.	z��~w(��`F�pZ�QØ����J^"��p�'���q��Gr��P񞆒�����_ߨ�|xN�?�X7��B������G�3nd��傪�v]E��pӧ;����/�i1�`f@y������k�D� �%��~;�̟Xy�#�L�)���!oQڷZ� û�S�{��ԉ������YVH��{x���s���%�� Ԗ�<�t{�M�3l٫y�`�1�ϩ�������޿��H\1��H��Oַv��K߹s���I\I]=��;�!��y��,��G���P�jfww�F^bD�
;��[��h��c�፟�7�8����II��ҥx}!� �a���������= E{s�Gع����!�%�U�p$(��ӵV��C\Az�6n(g����7�z��	�FNTa4�UO�m��:�ې}��7_�^�*m��y�9vߞ@H�=p�L�:�<vѣ�sɑ3�=���A���/��Ï9��QF���y ���g�G5,?����7笄D���f-�
���J��M͟���]	)6�߁f9E��(z�0�����Ĳ�����ӎ�~�)�������w�$�l�Z�n���*��G.��g�& M0�H���N��Ț�i�\~[�|Xē]+�  ����.z[���E�*� �����2ν�� ����֒�a��L�Z��B�2�
��@񱘽��A� O�X�y0����.t����v7��f����س<-�.�bB�wԶxʱM���G�\pY&�{�o�"k����ܼ.�:��v����}�p��u�3f�'^9�ץ�C��{�ee�����Ž�mjkvb�k#z�)���!V�M�a�z�@��0���g�gO	� >}�$�̄X�v�m�Y=8t�M���)�H���ʒ�բ�R�i@W�L������N�����3��i a�p�خ�$���v�yS�a���g�V�$Nr�+/w��=��N�5��m�B���+�B��O=N�yK�y��(L�K�M�/sB������a�++u���er�p۪<	oX��L��z�M��p��vXT�]�^�6G�~}0h����s�]�����>�ǌ�_��.�Vi4f�Z_��1�
��9n�-wb��錃���))2���ucܗ�
1��@�4y	2=H��G6�gp
���i	��7^glkw
���3��NV�n���ʤ�u�B�K��N����9Z#���g�KT�"��Pf)���A7Aޯ�=ASR��^`Y�M?L	0g��;|l�?�]x�`P��<�s�O$ ��gĀp�5]�e��`��ڼ~m�А"����E��#+}d�����ǘQ�z%��P\��r�U#L俕��bz���0D��/|�Ty
�}����������g&���f��S�+9��n���;اq�F85�Z�j�q:!Z����1�9��Z�;����{����6�Np$%ef�./wz��|�g})(����Щ e��=�`�G�v�����	3>N�f��^ġD����T�3T4�_�Rk� ��I_�զwt��"�?q(�:㌪P
A'� ��E�lS��z=��2i�k����a��P�
�y��!�^��PYw�Nj�bt���􎩩��@[b���e^�2�A��@�u3ͻ<�%�i��nLa'@0��������a���g(�`<	�.�o��:���d�׳�u$���4s��u�ͨ1s��T�:���ݻ{�F��;������>o�|��(�I�i�:EhYo�k������jo��p���z�4�a9��G���׎�z~L�5䍢*�6�?��X��a��m�uu���O�e�3h�0ve�M"+����:��>MSg��5x:�]��v!��{�n�x�����W�Tp�xlJ)�q�m��S��L)����wC�F +}��+�f���
�wh���s�k��9��`�6F��;(��.n#��=����C�	������`�j_�l0��:ES��h,$<�~�N#f��g�j��p0�+��O�T��c�e�nA��!F`�)r��l��Oc������{��ۋ^��^�8����KfFu����r���wy�v�e^�e�]R���(4|�m�E�ѷ��A5d��!9_z"X������X�y����ʓ��d/-�B3= &]�N�雯�}�n@�'���`QFTߩ[�Np�{�4 L��WL*��{���yrr�XJZ����Z���D��c���R��`b��W�'�?{.I�����7�~�ʉd��^��=5ϋ�Bn����x,?��m*@������M*5sqP�ʤ��a{0����S^y=�j�%�/�E���1V�տ�س���W�^]O-$�c��ߓЊ�x��q��<�ÿ��6�EH���+��r����I�sR\�����0�[c����N��ŋ|��{�j,�d,Ve!Wܭ�	B䈓T��c��w��o!
Zs�gE<O��T˔� ֓Sޙ�e%�i*�لvn��ǓiF������ r���䞗�at-�z	'9A��!��Ke9.ԡ׬<�A��wU���A��s7��V(C�+�Ǡ�%��OF�r�*��83Ѽ�H��XV�� N?WC��"U9	Ĳ�t�G�K��q�"-H3���s���E5�6���OB�SRR�	��ΐ��G{>  ��-6�=�Ù��Bm�Xz���z0fk�� �q����r�j�6��r�v< �2����Z�w�>@�b�WВ�侣a�R� �gFߦ�:��:%�5tz����|_��.,���K�F-�������i1�#33�"�d��-˿@���+�+�k��_g�}�_iW�sG��f+�v̿b6-�.��r[�S٦��ZAM��}L�(��6e����YJr��z�S��� A�����X)��먠��J]�cG���S}7�_��ŀ���T�!��������=ZV���ݱSSO�5h�Th��U�3�ÿZ��BM�f�N���������G�m��ۏӶ���;�n���7��&��+�P�Y<�f�B��N�����p:��<Bz���w�\Ȼ݃�9׃9I]a�T�)�-�0p���|+����+Z���D�QNV���}�?��#���te�u�A��g�,]�����p�`T��v�keت�~H��|�
65̮;@�:��g����zy����0B���V��Yˑϻ��O�k�<iwt��+�/3��חL�hٛd&st�E}����~<Pb���%%ig���t}��!���X�9��Rh��"ע���
��ChWy�����e;]�����nՔTzhw�֊�2^1�3�zj|ff��Ӂ�Y�����r)_�<�t,V�P��[�,Xj�qܘ-��TZ	�y��Ӝ��@�� �"���%P���>l����T��{�����z���+����Ӧ�gh���/Z<w�F������r]�Ph�=��b�U�zX����wƊ�N;ǣ��^�{%|4���s	�!�l
z*�� ,22��!�$�(�̖�_��%r�N�Aʿҍ8b����;�����5J������7ꧩ�NB�Hr�=8����Q��j<�ֿD[�,�C�,�u�6����./��D�:�UV��� �V��=���h�"V�����3�-�r�mA���h%HI4�	�����߅�3з���I�}tg��A+4������]�{�MCw��;�&��@�����S3[�O���W+eT=�����#���Z`��� ��V��a/4ڨyT����}h��2:�h��3:�m*a��ևV�}�q�F>��?�UQ�KN�f2�]�a�����{��֦h�ń=��J_��/��ս����$M�����N�J����\dP��<��������9���w'����h����<�W����3B�uXZx�c���2�m�Rr�~C����<,����ٗ��� �w��/��^*Y��e��8`�=-��n$���r��q�y��(g�� ��q��L:�����ۨY۳�A����Ʒ��y�k^��s��P��/~�>O�Ĵ�T����T�S�(y���En���>��xjy��nQ��h�5�� ,�KjF�$��'�!yڰ��P�*O=�79<�u���X%���@n6�{٦���UD�4Zx�C�����ا����_�<�u2b�ݯzh��+���3�Ә��Dz�1�s����ron���;����n�o�=��W[Q�l;??_{�Xǈ��7�	n�jZ��h��ڶ�T�P����6�=1þG_�u�"XY�l�`0z�!�������OwA�z�?&�:��2'_���b*�*�*�ga�zz��������"x\��H�I������cU���K]�͡8]*�!�|;�B5v�gp�2�3�nn����Qu%�Tnm{k�����J�)�H�
!�2g�<�SH(2e:%9��y�2%ӑ��<��M���w����u}_�*{�k=����������y��� �M��~���3L#��8�Gh�Ժ�^>u0��hyrU�W6ve����Lh�ڧ΋�2���$h���d���ƶ��F��y�V �.��XO�{L����y��������v������o�3D^y��{&�ڐݝ|D�7.�����?�{z�w��w��H���{��|�����4v�=��;���6+�S
��/�(�v���Q>��N*�2do_�7�O��REj;�g{��R�{:���nn������u �~܋��B��L�N���)ʹ�߿ӊ@=�[3_Ih@��czz�����6�j� �ȿ����x<EYl'n�3�n��8����|��J�ӣ��G��U���s7so%��X����@
�_-Y��c',������D�:��ܡ"MO�N���UCv�������8�%]��$zN�fS�M��0���:�8���q-����n���~_;ww��65���~_&JԶ��z[6>� ����?��M�*�K�&����D�Md��L�Ulkn?�k�Q*{ӌ���i�{��x���{'i��)y]�HZ��b���ʱ$���G�~;��l��:@�;;��5ǘ�d"�� �2۾(�̰A� 4_n��*�>i�{�e�<���.V���KS�c��I�����"V�=<�G��LĮ���ԇk��DT�����@f#���k��Ag��x��aMu�^�ou�E���qt`�O����=�=��:/E�����~sx��P��yapԗͨF��`c֧x��?F'x�>ǿln����g)�\([�~z�馨����-�LL'^G�x�+��{+ȯ�]��.�z4��,�]|gI��H؏#�AD)�u��-<�凩a��w���8P#�C�p,���|�p%�!޸@;!7V����.�T�ǡҝ<��_�%��z�/��j�'n�:�K�c�G	��gc�_�0�u�4�]xŹy�C����[s����Sz�Oz��%N#���#��G�W=�|�*���^t-���=f�s��(��`f����/�{�����(w��Vδ`hM�'xC\�ja>{n�nW'� B���=�7��J/Ǿ�a��&߲?E�c�������V)���5��KY&�Uӎ�#�gy����EK���^��xL����sT�Ǔ=��E��ru���DP��)m#��f�#F�	=�����i����%y(g*x�o\<`j��j���F���F!�+��>����d>
�f��
}#�Ī�������E^����\.�a�980H=C�P�=zf�%po=�D������G�mvڄ�f��ٲ��!Ҥ�ݝ	<�U���~��2�0�%3����L��d�wk�^n�炷��
��9����z(O������ �����{�K7D�V��[o��s���/+�U�����P�u[	o�X��m�#�-5d�%�yz�,5Vi#PE&�M.���f�**|"��E�"��3t�����o<L���pX]i	�Gɀ��F�×��|��|���</�P�FJS�R���G��?�Pz���kl����޻�{����kY�@ݏK�� ��Qij�CK�3��%R!��w����,=�ZYɃ�$ɓ�۷@CDL�~�[�pt�b[����)m3v��o|�Z9Ϻ�7��������踙[Z�r���@E���2��{�k��Eh��z�V�]C���PWgJ�6��[Vw6��E>��8sP�P���h�	�x��[*�O��v�cc��z'S��@���Vs��~:�@�5u��'Yrx�拨��l�_��?�ڽ�nq��("L؉qV�m� ��{�(x�2��c��N�����6��ǻ:G~���?O[`\�����]��7������T͔��)���8�m�Q��(
ն�,G�s�Y�R�A/��p�FaR|��p'����;��٨��{`ew'M���&c�u������e %�ݍ88Л���r�x��)��������G�]��4|��,:d�zRh@iK�ݍ]��c.q$#1�Nr��as�d�fJ�v��Xo�h3�)l��Eb����q��B�_S�]]#��S�����#_���E�����	0Ϳ'n�4Yꋡ�����ϰ�FOj�o����W��8�4۪k�is(���7YH�v�e�?a1ů�R��+o1��<����Y �{---�}}Ǣ��8�TN 8^ZG�ot�I�	�����g��0���M26���24��I�K�h���g�t��P��)�Q���Dﬞr\���or8��5��F�l�j�9^��y1�k�=&)Rn�z�hʶ�ҏZ7��(*�y���"Q�}H�'�2�/�I�DI��y��6�=�Ex��9�C���QZd�qzl�MFq3�t��-c�E���)9�hn��6��*�-7���j���'��I��
(/Q}*V�����,�8�����""D
^�����%}�ZdV�%��5/�J�T���ÄV��*�	�ҔgMMM^,�bt[�� ���L��CHՠ������V�@n��2��Bw�<����
N(��X<|O�9.����Sa*���|2뒀����thۑpYa���8����:��tN�XZ^�$�Dע�!67]�h�*d2�X��5�-�{��QG$͖
��7�3�uD#�`��p�9Ξy��'��@{[[++k�쬈В� c�r���g���l��X�����i��ƥB
n�1����Li+-��8�(Q����-N�CC0(gi�f=�1A`���Ĕ���F-�{z�}D v ��a�m�� �LK����fs%��=��h���*�W�������Ъ�y�t�r��`�1ћN�}�fe=AD�m��Ԗ	$�+E꿃+���
QI䂹|�� !�>�|:7m�]̺{M��$�aU՛�v���z��[�9RI��ݝ�s��uw������/e�����������b�p<���J�)��" �|��φ7P���<U�ځm�������,7�!q�/#m�Y+�-$����rk}�n�ĩ�����?�t;|8����. d�	ֶHl�H�v"3#�~Jӧ��fvu���O�����Ig#��4�ݪ�N�j�g�Тk�[�L3	�� �8����Nqq�}���(c\n�����잨!��:���h�}�d�O�#��ш�d@^]�q2�U�y�0=9���kL뉟_� ���qn��ǺWw|��N�C�>hV���Y%�+�ɼ	�h���>+����p>�:�R����jѝ�A�|�^���bIv�,=�ZL[���~�z��W9/��p���	��B����T������?{��� � ;n�n{0�y�F�&L>�QDvm��҄8A?�*[�̗6��������Uc�5؏"6-:�-���V�I*�G']�AV�8�G�;=;�Oo��zf��y�P�N�q��6���������v��4���$C�v��3*ɏ��af�#_�V����k���2Q����_V�)�QNJE��GB����;F�L��4�ۙ������nݕ���FC�g/����r"v�k��l���39�����S�ȯ�����q]��g ����e[ngh߂b�NbH�d|�A���S�U�'"g*��#�.�#�����lO�:��y�=3/�#���.�41ISK�Kp�"�O�1L��m%��F����(>Z�9���E�NNN�<��|��ѵ� <��!W��̨{	���;�V����	�t���*�s]�8����r"�z�n�}+6����	��`$[����S���W�����%?�_sA�Ho�+{�R\��tZ�˖1n$�<�����π)�U�#�����@:��ȁ�j�cu��Һɷ,s�����Cј�])��I�lT�Z�9F�s��N3�P~~��9~��⁵�L�L~�=YU�)� ����?w����Δpխ��	1�"vB�!���������O��r1�:v�1�#�Gښ)�H�NO�lc|@�d�ܯE��g���K�"���A\-� ��Skto��g<��^�}����|��/sVZ��g�߿�����fV�V����ąȩ���������_c�N3d�	v\���L��Pі4��ΠS�t+�Q���#�3~|�Գq���uAn�$�f�:w�vJSHl,{fnn��S����S���eh��h�^�M2;�^�OhLr��hw������>e1gSs�T���=4����Z�F���7�г�9�inZ���i+yhL·�+2����I���
��lX��م�s���w��)��R��H|����p�ʂ��S@���z��gH��^�W2۾�6p��Gi������CA��κu�N*�ܭQe,g/	2���4ƥ�f��o�Ϲb'a��@Z.�8��N�/
�4P�W��9�illl_Iɓ�&�����$�NJ��'�����/
./,�Q�;As'5f����uX��t��I�/7l|��y�*��qB�C���(���񔮔<�&U9��U��t�y�vᲛ��eYjn%)&�ra�	��v�fP���!o��W�O�m�f~.��~���8��I����m�����)���z���C�:W#25���$Xe0c��D�����Pw��D��������gZ�Q�l9=�}&����w,��V��5o%�b���n���e�<Y5�?ZQ5dR%=�a��zN=��+ �GM��=����Q���sn�ٷ3\�=6yH�Sx��s��h���d�.�F�ß��a[�fI�x�Szݍꨠܻ���1sHռi��ƴ�S��]-(�A;	�4p��g�Ϳ6���my~�L�Ӄ� ��|ȗ��ӖO�%L�ݽꡯ ��C��>(���y&j�5���Zzh���FK�^���zMII���^�e��e:���7�98>)&�SS<�����XQ�&1P��w`�	C�*��L��$DHd���k�tήT<�"c	IS�6tus�!O�]���EM��ots{"Qot*8�u�n���tW���8����9l4���Gw}�LI6��Ie�\�7ꇘ��)'5�z ��|=D�����>]jp\2��+��4���>��t�ʟ~���*t�{��
������}#�3�d
�Q��lPV��V)�:�-�S�M����-��U��_��o7f��|9�f�9�,MJ%�R�l�/���rb�&�xv�T��Pe]�CHf���z�)����]n爾�P��C����I�(��(�"���"dK��Yr�W\�gf�7M8�&�Bȼד�DJX�z.�·���z�<����e;ry*J��L�f�i;�4�so��fi�9���a���hW��ӕ��ŉ��+G@+8���1��f	��%��WGM�J���s�?�	ypF"�kw��1y*ͽ���ٶi�k|'�,�A�a�����m�-51'�KD�ڍ �ʏ�Γ�؁����L^����k���0���.�7pi�q������d(��>{ۮ�#�~l�t; ��xh�P(m��q��+��Y@P��#0'�p�>�%�5�f-h�:���+쉨�>�4�X"E,8�\c���\f?NA�z#N��o�Ҡuwpv�<\��I�C����ױ�{�Bs�h6��o��e��C��ɷ�G���ft[V��:��E
�oQZh�w��F�S�[
��#b8c&�{����Z��S��Aw+�.|@�P�]j�[dAV\� �y?��GZ�S����&�ZQ�x>��3D��U�=��=�� �����j2����>p9Z%�\��p0�<K#��S!eeb�;&�AU�s@�rk�ro������_*i���o�i/�[�C�S��n�kY��݆�	R���=�-�H�>b��"[�n��Z�T��.ۚn���&4ƣڪs����C����z\��Et__l+�z�Ll�w1P�PE ����޻o�@82 �EK�@� 57��M��]<p�P���n��c�ج#��<��� Z��2|�Z3�\P[ppp9i�K����hh]��@/r'Nw�wJ�x��A�����h%쐩�)v��pK�� �*��gf_��f:]�{!ߚAj��gW0�X a}2�L����=-�)����������d�k�_i>���};���u"���ENNfx���d�A,���Q���ޜ�u^�@OdL���g�F>R�<���s�ι:)�1�F1ei:76\�^>pa��Gwqt��훯%�e��&�n8	��Q/��awF>���w�k���r�

��C��a�ٖ��膔��v�$�t�aF|��Ds����tg��˘�Nn�Ԑ�6HCg�_���In?�s	��L\�H�D �r�ne����k�+..P:�R�ۤz�x��_((��h'��Kl�eb�]TP�L�
����+X�S�Z�W/8J��:uA��V6�\$d��Sk��x�5Q#�/(�-]\���:J������L�!^-�0ǟ�
�v�|F�,I�i��v���⪍8��@�3Q5��NwŠv�M�f�1��9�V�R���� �~i�ɹ��YU)G�u�n�U�uvg�_E��tS��"O�w̥a�f"�PK:Zu�L�` ���^��Ք&�Itg���o�'��%B��Nkc7(n� {tq��V�o��8u �\��w���.����S���O��u0C���&Sg[�5���o}��p�Q��!�]�6�B��kS�;���S����\W��%����񬉉�tA��7�d�z��O�Z-�Ln).rG�I��BTO��^�SI��9n�/z1�k�(�M75���;�>��q�G�`ZV�9���^m;t���N���Jc|��y�%q��M��ih����*�b�7:I�{��|40@��Q#�g�
v�?��$`-���5�ӠI�{��&	��n����V�>��5P؃�0��0aƨ�3@CYHbb"�'}I�=�<��WC��pF�����.9C���tcA�}.N-�|^����>�		��lb��rv�	c%��3L痥oH�jvU�6�}��i�+�kǨ��l��O,�Go���>JCx<���8���g��ɼl:�z@7{��g��o����9Ҡ�+�Ɉ߫s>��aI��(yϴg{��}\���I'���N�ԋ�c���N�>��B��h����	�5̈ܬal���zt�����n�����j^�:![�$�.����l�����������ch��)m�b�I���Xkʰ5�1�����E��A��^Bb�o��|��B��y��&];2��|<P��9�}�N
��0?��;2�������8Փ�� ��� ��%������U��O����e����i�=?b4��\���^�S�=���<v�3��kf�\����JbTvS�v���T<��� c*^"������r�$��-`�u��K�+13��k߱@�� ́T@�$c�\�(mMS=�-WOmϳ�גϣ�$&1f�A��?��ްtT�e~�x+:.>�4�a��,7|}�g�JCڄ�!�%#��Hbr��
��U+�r}�G@9Gǂ�4� xm�h���:���̌�������}��Q����Vm�Y]3yX����3�X���|�}{^��\MILm	[ݾ��5%zn�i�o��}��ܵ�RX�ufGA(���H����5��!�`�x��=��[,���d�ch�"�� ��wY�� �)�/��yM��2��Y���_s+�H:��vؔ]SS�|�8ݙ��e�|i��Eʗ�̛Xl;W�[�����Պ����h+'%'�i�ńi���rVL��%���6�`>{�l���y)���������e�/"I�c�,��G���������l9�A�=a����n�r���{���3�1I�$I=�P�����-H~�ƣ���i03�s����F�-��=)M�z���p���4���(��S����˩����j�4}��"q�_Ces�����PD�����gdC4�۝צ��D�%�+�G����/�3��E�
T5��<c�?�����P_&�Y�	����M�F���
z�������Ӹv���I��� ����2t�c���>k�\Nh��1)�CW���r������ 	=7� z8�������~p�����WB�Ys�۬��,2.�>��$TA�xB���������[�$#GGG}�"m�D�h�LEŚ��*��1_�E���[Rc���3�c���_�6}n0}0d'AT�(�WSCѮ�0�p�q�48����nb�NN����ʆVV����z�S4S��?�{�R� �斏 �L�å����k��==� �x��z������q�a��r/Z�Oƪ�����lm��m��tt<��2q'��O��8	m�`b�F���{���K{Q�A2�{(S=���
�m/a�&43o����o9��N��]��#��w'2�P!�[.�c���mȗN�"���߿���!\�k������r{�����+��T�q�݁�I� �n2��>3���|�����g�lo��>V,}x�T�\���|�\��5#c��&&�q�	n�x��JFC
����D�������|�]�z��(,,���dΧ�!�u��\^�o�Xm�1�a��s�@FiǍSa�"�Pm�R�[̖KA��uuu]�ip�=�f	�MD� z����r�M�<|������q;.쯨�XklkLʄQ��/,���ǭB��벂>�����V�<����/ ���Yۖ��Ⱦ�K>}+¦��"̴sq�*��}K3�%S'���͛i߶μ���"/uX'tL���C�O��_0�J�xF M�ͤ�a�ޡ���̶���ãy��B{;::�ʴt��&㫉�U��]�]��K��3�w��}��]�L�R�ڧ"�����4y���C�@����1d;���x<��P��h�b}��9��A����5Q�5Qg��$���099��ߥ��]7�a�{�X�8(v��޻�;�F���]�J��ܨ�r,��*�Z������������{��Ԅ�#ɿ7��Xa�y�%� �q\9䟖	D�����s-�͛.�i�v�E��o3��R�~:�}�==T�ɓ'�W�+��s��x�Q�V�lʜF5���O�3��<��
���N��&�BuM��[h����?ۋ^���+6uw�V������p���@%��?�'5ȫr%d�i+��/##�a�d�ˆ�N0B)�����5��!�P�{Z}�ZC�]N���H��y&+��~�	��?~D�rr[�{�N�rj �����Zc�������d���� L#���(��m~�/久pg��[��NCR�����Y��B���)�o�t�v�1��)����6��+%�2�!�Z&���(\SU}��*�h���";��V���������t?� ���� p�Z���.^?���"��fzv�ET'LL�˹��:q����,����w��}��޷��<K�ΤjNhy�gh�]&���iD���FT:���e//��(�#lx�e����������񱱵?��Cq�;V�=~���H�p8�	�Tf�C����'l��rܗ�@&j�Ͼ(7�nĉ?��P*q�`��#dP$095u9�I��;}�G3{��Q{��y�m`H�KdH�`��>�W�xC�����s(�ٗ'l�
(G2c���\��Y7uw�c����RG��a�&��b��fP��+y�	���="22����M����X�{�M��8���B��{FG�|�}�P�zWw�0��r�7j{��J8�Vl{����HK��qqA��ښ�A�q3��0ZXXd|�r ),x��#�_
����b�R(r�l(I ���<���(����Z(��ʍ�Ok��ځr�]=�v�������υ�m��~��"`@b���{���Ǌ�����O��dFEEEFEU�/������C����X����I���K����L�����3*w�g��~dh�%K���J�:9���� �n�'���ė�z�BS1�	-F�wn}<هF�o�J�w������y�D3��{����?�9
_���vO��[Yc����3i/�kjT�QB�'8"�ۛ�"_�:�o�݁��$���&T�YH��/X�"���}o'3����a��
��`9CN�Tӝ��+�����_�����z����;d Rhi) $`��%�����˂���[�w�+����V��sUm����4��aی��W9kr}c��^M9�:����D�L�w�dn%j��AB,��BR ?�q���|4C~�6Z�0��̀�"^�f����Bo���`*jhn~
t!z��������U( ����O:םo�&5�q��v[�P�,��k� '�żc�4������Cn��ܫ���#��Jѷ��� i�g³��ӕ�Ӄ~*n�ɑId�S�\�ʽ����$W��_��zyOETC�ж'@)Fp�r�I�99���n{ �h�Gf��Utm���C�ܢ,��>��q�o�w���/��綳)픟68��n��Lv>�,8x09�@%0��TM~�*�"4�����k�w����-=*O��d���b��+�L�7�����ݖ&G���}�I��H�Z����9��Z�=�hoh�����=�~r\�?�C�1}�
�w����X���44,���;�1[�	�C�|n	�H0䒪�j��5�D����Ba*�[�[&H����.�;w�P��j����菪QDN�t���' ��އ�
`�U>~����O=:9Ay �����ւ����ԌJa�m����F�X�*������udW	��
V�{���kjk/��չ������΂ܱn'vY��MEDaڂ#�a #߾}QEd�,m�Un=�|�pm��f���;�#�^olieU������e`���>��"𳧻Q4P3eQeazo:��Lŧ��Q�Uh!�����_�J���ijialIu���f5�X��6[	�}�1�m�6.(��&0Y<��8��v(�
�-����H�G�vvgP���N��tg��l*��clsI冨��v�.�ѯ���.K4�622�
����e�c��!//��g�anO���j7277�Wx�� ��_���ѣӌ���&�P&�Q�8����X��l:4t`R�4ac���b��̤��;�������V�l���������W�T�Ԇev㺡)�G=vVV8m�L�9��F�xy���ϰM�u��RXϵ��so�dl4��M�W�>�s$#�0^���I<5�q�z���_��Y)���̶��m7g73ڐ����9[�ƙc�Gp<���_�����xH�p\�'�
q��7~�JH)7!��^E�f�C�����Z_c�5���A&Ofֿ�!v2�yV�DCp�)�?O�~ѵ2�0�2�K���'G�^���2A?U	��b�A��qT	�	����ge�C�-�<���h�,�	  ..��Ǆֻ�q3�a�C7jdi�++ܣ�q�<�_Q����3��,�������L�e��l�P��i�z����8_D�#���Zc�YWk�8�:\P�F�!p�	��#%n�)ɇp����uu�0C`�FΌ2o;Վ�N����|k�>��jZ �B-0(㔣�H"�\dɱ}
�rc��(����	D@��n�N�\7���ŉh��@��r_���;oУU��Vwǔ��${D7�7�	H+�RKOuUJ����CΓ����R@�|q:�<Ɨ���ٖb�9�7�g���QZ~@)��L��;��X�u�`�v@睝�'��A����������mmo��E���p�b���:�+cI���,���f�\p�T̌~v~���J	b�Y?���6�� ��T��Q�6�k��[#�h��7���wy�
F ���@��t`�s<�]!�P�@1���]�.p�6��;��͗܎S�D�r�ރ����h�H'~������������u������A��+��E�y������v�*���@{�e�����LS�裞`��Lu55�D�*7F\����"=���]C����ԗ�����]|9�%�?���7*��ª�½D"A��ރN�Q�H݆z
3�O��,�Dp݁c�\���+��U�(���P�g��1ۤePƯ��	�{�bi6�N�(,H>��J��f+?�H}��!�9�p�=Ϗ���j$�l�2�_�f����:P7��\�܆4������B�����d�1סe �:LhaoMo$/�P����>�������$��u?�!�zp���p;�H�%�6
�T\Iu"��皙jizm��Tn�j�[qb���j{�V�.b#������~�-w�s�j��
������w�9�#�E�]@˵ƍ�;���s�T�R?t�c��Z=(��]L��{����@HPS�?�xa�n%� X�ݖ�;s65��&&&f熪�ra+7R�3lM�v�E��;�(ή���%5�>sƑ�+**��[|��
��pjh�1۪���� ZgQ�ƾ����rp��3��x6K����f����x�	K�� S�1`���-�Tէ}ɯ؏SP@�m���l8������^иQ�-�"���R�$QD��2XnUO/��USZ�Oȸ.������#����E�(��[�`ڨ�P>��>-F�Ipxd$��*x?n�����Y�ZS�[��$/�y�w<k�+ww��a�?xQ ��(�_�L�w�^��}@���{	�mjjB"��<����Y�ڪ��>i��`�-���s7��:4#v��Q�#.O����ʈ��1O��#�R�b���$�痢����k��o�b�$P�m� �o����`)5�̈������_rs��Yw/�?��"�T�sM���x'����������Ւj"x�_��4Μυ�X�O���v�e�4���:8�C�A`�l��F�쁔��trk�����Dzz���0�z�E��/�.��rC�"	z�=������ &T�y;��_��P���:�����e\�����,N��n���SpEK�8Y���$�����.���3s+����K��"48_]3؋?~|Fj�Q	f_\��$�B�D��;ղ���<�YK?��aF��Q��&�=�j�bI�t/��;(À�'���տJ,�V���
y�A�s����������N���0�\=JS|(wը��s9r�F�'Tt���6��gDΟgDN(\(�:Ѝ4���ލ}/�箢"���ڀ��V
g#P���9E}�>�=�s�����>�b_i����ϯ`8���/��ˌ���`�)�w!�j���إS
��1�UL�#Kf��nt���e@CL�0;�F�)W�E9)TC����}���Cc-8��ڋ���tJŪ���(��;7��ӛ����'�<T�Y�Բ��&���*�xΈ��
�1������A�fR]�{�� ,lܳ�wu249f��.�[p�vе��$�ɬ�k��n��)p]ktZ���m�!����h]��YI��ט}s��,�2�8�7�Y��MKR�R�]�n�r��V�Hs�@��=�H3E�h.��L��><�f���[\�|�-A �y��,���q/�sf$��~�Mξ>M���P2�'М�����������y�b��C�[��^]��w�K��s�$�_��2Ϗ�ͬomp�.�z���2��3�겓��k���=�����A,m��~-���W�Fxp�J-h+�1�����I)hA�赁�X���<�F��x��ɓ�it�i��s�x��l�?H��(�U���̝��+��������8��tv
�l)���X��}�_tr�7O�qq�ؖ����A��4��8���q��o����׾�#�s��k6�L�=�f���	��x���h,;]hG�Z��eu�Pey S�fJ���$�%?�Z�b���1���2����~��Pn��t��Uk�@J���X:Nž��/��Jk-�]��~̬�՞k��a���o���=^`�-M�`DC�h���*�G�ҽ�'Fߢ�w���K%�Ŷ��Gvj!�O�ǣ��S
��m�0�`�@�	�}�Ik�ϗ��)EK���n�e��^܌.�!�
0� ��d�$��/��<����#��#�JI���������D�.0vh}�9#��I\o�AD�ꦒ'�YS�@�7��gQ_� ��.@�~D=n?�������J�~��x�,G5
���A~	��H�U
L�ag��!m��"q�,�+fh��	�9��A6�ve��ϟ?+�?�^[D�Q�����2�8�t�_+M�P?������m�2�j�E�G@e�:�#�e��h��y�l�,"r���S�0�M}��3b�")�D�Y��S�Fk�h�պ��IB���U@?�o?�.�5�m�k�+�P?���k��lђV����m�/ZΠ�w&m9��f�o2Ƕ�ű��/�E���D�w�Z�R�ȪS��z>�|t�.��6ې���C�|�)��5Qg�Rff&�@##ٻ���U�{s&4� 0�(�1��r(N΋#::}�5��O���C��ѡMkd�����Hٔa����CD�oHP�K��H����ƊVJ:����]�	BNS|V+�����k&12n瑯��AB5��@Ã~����z�n����z�qf�rvى�L���"���y[��rdll t"��7� ��6c��323C��G/3��8��{�~�֕�Z���J	~����9��O3�S���Ͽ��m��X�m7ڃ��X�G�̱R�G��v\�\>C�@#P^^>JZŠ$��k��\�Xa�)}�T�58ྈf�d+떖���\��f�V��$@l�KW���G��hI>|#�֟�
 �8��=VD�Bۍ�a�g͔�^�1��(�m����/�oa�m�m��l����yQr�	�t�6�~?�n$:��&^��O�}�	l�����:Ց���%XJ3^A���30,�iR��	fv�Zܽס!�((`��P�)��>�����$�^k�h5�b�C�����!`����mv�8z��TP2�C��8R ^W>��e3��*T��4�鯖��魅����S����)K��(�^��P�L���Fd���Y���[���Ds��L/���.M���a� �񒠽++t#�N1�%��>Y�d�V��@�T��eV��p7��nʦ���O�_���k[��� &�~9ʀ\?�*�W�(I'���H�~�/�����A��.��xl�bѫ}�6�^��9��h����u%�a8ۺ'h}��kVؘ�s�E%����A3e3J� Yt�ћ�E܀�z�1U�V��8e_"�`@��� �K	��_%Q5rU�^��	}+Rq��y�@(�-:'��bdY���R�fZC$�F�̃�WzS����� ;$��J���*��Fo���ۊ�fMD���P��OaO4tqȺ3C�QtF>���m?����� )��2�
T��n�%X�R�@�3�8�Z�hY���.�ʹ9;�B�Pq�7�3��9�w������U�^wcT_0bs�l7���PY�o�ƚ��:,��I�(��D����K����Ef���O��{"V���gB���l�؋$z��A�О$t�E���f���*o�( *��&��I�7&r(���8�����J��`���������4|9��?%׉�+�~*P��9;X�6�ѭ�pi#ss�Q셠k����#2�};t�Q(z4!��J7#�@_�/���Ӵ��p�?
�.�����u6JNk������ �y�	���ի�ɽ/aw��G�"�{<Y���1a���WL�G{��+vgZe�������*�o�3|���k/�3�h��&A�2D�Ñ�l[�����$��WE����Awp˸B�[�<˅v��­,����<Q@�.$�p�6�IB����"���0|��,8w&4	<��<£��0���K��X��c���B�Q]�sz������q@#��L;�� N�T��1T�pc���h&���0�$��lZYg�ޭ���0@���`T������+�X���D�}`n�����/(7ZD}<���nT��X��vF�$��&?~,O}�7����7�T�d���ޗN]k����k˓����ԫI@J�� ���@�1���	� t�
y ��cok�o�4Q���G3�7ʺ��ܤ��V���w%�i9�'��QF����KCW���Ǉa�d��D۔!�w�7��wJ�/<�^щ�ζd����E�m,�6
��7F=7髦��b���@܅**1�R�Ƹ��e�����c��J��@UC�R&~�rS���n��]Y&l_�C��]Bve4�� �#o �`>�l��š��03c3�&��MD/�244�ZQޗ�����
�I�Q����-~�,Z�C>4������]��BVt���uh�04h�r�N���N�S����!��?@C��+�;�����+r��J��\؎�J&���B:��h0�`Nǣ�����9�M�DΝ;�%�W�,�2�%��X�wb1����<қ���`T)`�]]u0D^���A������$�[���f,��(O��J*ڃޔ�;��ʊ��� �Q�p�n��ܠ2��`x0�)�)r�,r.�&�nA� ��ab+m�.vL��;�h�sZZ�NN�-iwΚ��B/É����5��U�q�jx1J _FGb��т	�e�㑿�7�~�߈c��E,��;���}�N	PTTT��Z�_t�Ooj��^2֙<sF�5�e�L�L2��ENs;��pw�����ԣ(��--��{�7�q`"E�W�Y�r��!�;	�(*��r���HW����זa���0VD9γ��@���ѱN�����]�P�c���[��W�-`^�?A��g']���<r>�𨪺�^,���`��uP��A(�+7?�È����0��ê��q!�F���p-iU��̒g���A�y��`WQK��)�� -�|��~]\�c>;"Yp�l8ۙOh��;(�<"��Zo�8L^4��������De� #���Zl�6~@�� �hϣ������vN�J ���3�����4�a�xs��D��(�`��g�~ʭ�*	%,V���y�&��<T`�ѮP||0R�T� ԇb�x�=HII�mH�������*�u ��Elha�th��sPST�P���E���8:u�E��Y��aT�F]H=��^o� ��ާ��;?���N�y_JkAC[ h�?��gKvr�u��0��c
<��؟?fAܘz}(h�8Zio�2��)`.А��;g� T���H͡eD+ШD�齂N\�0@�"� �E�:��U)�.H3R���D�����56�\P��g6&�����V?�ۢ�w�@⌌�C��P ÇH�-�8�Ld�R�6F4S�?��ox����p�����f�kc����������C�2)�@=r�+�y��䵏�S��r׊o�4�����wc�Eߟ�*�v� ����՛�eM}}O����'[�Y/�0�������&s����E/Ʊ��VF˷`��������y&/�E�UX�NLL��S�ȿuj=>�w���Y~�Yu�K��f�q���\[_���EA����݅JU�NE^qN-i�Ҋ����Ȳ:���H�6�'j��RYzb7w��cL������宋�.l����ω��dZ��c�U����ʻ������wf�����!��n�[I^9M�w?}��t��^_��5����z�Ћ8H����f�ݻGxV�YV������..���iسaǰӭ��챇_o8�x����b�O��ʵި$>}l������)�%�߰I9���fǤ�{�=��r�(�X��M..N���^����)�RA�;v�8?8�/���߷�ޢs�oA)�}���)�,����.\u�+��pt\�Q�����l��_�Uq�'"�ٓ���)�"�(�7�'�/�Vl�֍�����
febd����ڊ\��7�p���#�z�W�n�J�[j�0Xɭ��&�fc]��j�pqƆ����!�{KKK���d�|�2s�P_���΋s���055}(�޷�G.lp���ؽX�4�䩃��500��f��N�>��ꡎ��5��_�]f���~mT�8|p~�Zr��C�������o�/�b{0�I��>G�k�0-g7�#:+���U�D�J��!����GF}�ju��ċ��u���v�����kF����n�Q�_2�\��&����␫�i��:9������MHI��Z�r��0p�j_��Ծ+v76;���{���Ij��g��W�����$O���5��
ꩬ�W� ��u�
P/�]�
�c���"�������o~k��K��n�-�$����o���D����t����Ф���&�,��a:xa��ę��%O~�'�`ns�~��~X�aF���	*p�Jb��nLn���SV������&:Y-�A��A�z��m������ݝ;wVF���i_���Ż�/wn��'�:��7��')o{��R�Ͱ�:�ô��e�]ң
7�|9)�z��8ne}.A��؅�&�<;�X_��vd�j��~Z�X��ߺ7�w{��������~���#R� �T��E��/�`����X����T0��C��{�����϶Q�7�Z����	���|b�TZ��O�f+�!��Ɨ�eb!�?�/N��xZ蹯����4��컰ї�������

M�#�,�D��Vo\7�\6���Zy)��m#�M{����ڇ.{���;�Su9��u�7�N����������[3���&>�LX�v[Cߏ�z^��S\l�SU0b����`�l�'�͐/H�	yԣ�,..�N��b���gJ�9Q�qA�֒�t�J����=A���o�]�{P���;�(��xM�ל�����QgM��>���5�?񝸀���##1L���v�Pr$v�+l���a�R,��4��-�������S����7�U�$]�9{��go�c�j*u��n�؋�<1����K�����P*�9��H�ߏG��j1�/@ڜN(��8�q@�@~R�W����������r��^S���P������?1�
��&��2X�8۽��vo�ݔ�l�F����ʇ.�T��s�e������k���7�����-
�F\s��֟�Cپo��3���^KHM�R�(�e�P	�$eˮ�죒�V������I�b,%$k	S��l��3���������yK����<��~�y�w����ҫ,�_s����^_�4�G���#徱�O��'ﲾ�K�!Mx�"��߷�D7En����o�ѐ�*�1P���@�*Qݎ��"��Y�D�X-M/�t� =�ssPY����\��������XO���_r�N���T��,�iv�<�P{.j��CO�����0�����6�y����6������a%��TMi����n�+��!Bp�ul`e[���Gn#�ߐ�_	tq|/�0/��6�yA@���?t����k�v,�� �쭭�t�{c��A'h���+�����b7�w*x74<�M��7&��dR���)����%Z�d���Ϙ	��P�+��}RM	�G~TVv�먮�Aݎ��K"�J��UG
ۏ`s#�6Ľ���;�=��_Hޟ�`f��|K�������2��bB���hpc2�19�HA@@@��� �K���L�K���c�	q�}��P��W*��9`�Rw�Pn
��������^X��꿳�[��UZ�#�3��"=�~ȧv��A﫡�oߊ-S<������~Wv�-�<��G*I?��n:$'���lUSs�O"��۳����1|Ev�O���mZ:�,�1��C�&z8�Ŗ��'���7����'b����(Q��7,g��+x̳t�]��`pc�U������{S���ް6M,'�/,dx3�P�sb�N���"вRP��`�]7���m�[�e��LhL�(��WN�	���1����+߼=�]��JVH�V�Y7'�����_}kpC�7����6rk�	��1ֻ����'�	�+\C�>\����L�	j��DM�s�����
��a�꟔�4���8Fs1A"�ߒRx�R!�_�~X.7<��iV����(Xyw�@�t:�R����r�M�����Muԏ�J~Ք΃����ׄİvC���t9v����Qq?�_��
ݒ�9TGp�tl����oB�X?��'+=�����(���^�>�����aF����+\���ka��b�;�o����֖�"�ʎ�X��{]T��^�'_Pn�7���/xa��r�]��%Z�iiK�;n�	p��mݺ��0~➭ U�'0L}{��y�,�İ��������U�|�cN������xZ�Y%A\��e��&�:f�#�`�|�ɯ`3=�Buը���?�GJ�U��xA�u+���J��@M���V�������T���U��!]�����Smh�`x%,��K�}���|�R�V�v�nk���yp��U"���n��肕�g�AJe�l�����*��}o��g�����Ư��g���Tr��'�A�.�'�5Q�9�[v��ښ���O�=�����=�v�y2�7�]R�sq�L7�1�J<�,���$WK���������Pm��9��1ڦ�^�9F&�����:�j�!�J����m�;����Q���+vVK�<�Z�p?Vf�������t��.��i�5dd��s�-��Haͺzz�BBBv�H[S��K嬕�nf,��_���{)BdGGG��ؘ_A���D�_y\~���s��cK���T��X&DvZnL	t#vq�|��dhXX.Wx$���3��������t?��������1ע�����l����8Ḱ������)��8�s����j�5���
�Z�3	A�ao�#�K��QCb �(�k�94E���X�7��-]�Q�+��բ�JQ�~�ѓ�H�׭t�6bC�s.���c���Գ���-�(-���J6����d��1#X2&8z����.ثn�Å�d=�>h��&��zN_M|�����P^̡���")n�����2�x�pՄ�!�ګۆ󩪩҉.��3����7��F���(�y)�͘1t\�c�I���S�|�qq<q		�Z�BZ��ҽ׭�/��G���i�v���	7К�0e%%_Q׃/B���>�l���=p��jFUD�݌�Us�|��+�����_:�I���X�M�^�\:����	���ַ�]���#��`(�֐�r���{�/�e���T�k�ช>ܸ�K	|.���۾�^�KD\��m���=A��)���������7ov�֏�L���?�aR�!��\���h��R���Z[���D��ڠ�4r�=��m ��אj��xUY�O��![76����B�p�෗�gf�ǓVl������8��e�ܞ����X���:\ʙc��
�+w�|�{x,5��9�J�
���֞@yH1ݣ��x��A'.�Wܷ7�j��� ����d�����5e@��^��~��@\����[&�]�x��4�V˯�9�!2Yvq�����v�Ct;��`�&�m���H-�������W+���988���/�k�ψJ{�.T��6\����K$��i�m����#mgl�5#+���<��iR���c`��)\Q��M�~�2r����s�߿;��߉�8ߩ�e[b�Sʂ�6P{���Gy��a�Nrck�ث�i���	�۶@�K����u�D�T�d�c�� /�d����?��4W9�3�F��
o��~�{\���N$��p<%Ҡs����9UGUl���[`�oC�	�^�x����x�ӃƻKI�KI��k�t@�F��
����>���?�F��u;�D5��fS'��"�G��Q�=M>q�zFi[&i̤��wG���w7���RO�T�*�P_��-�-R�|�d J8G;�y�P�ap�}��;�e�Fz��J����H44��=U������ �`'� !]��t�:V�-��Pd�j0�]���tc�2)�Mc����t��(����x�P���@��>��vF2?�0�z�G:}si$&�3�z{x���J�h��	 Ѐ)�Y�߷)���}�
)�NwM�UPZ�R�i-_����~	�dm�VGQk�C�waW�������B~K�uV�=��Z�Ýy��a�sn	8��-��v��(�?fV9d�4�K��wn��	��џ�yk���_��76�Ⱒ:�A�3���ONr��Z
|L��a��`���>�c����jMąƻ�b��+t�U�0=w��yߍ�4�)�n���v(�M���/C��{��#A����W���`Ej�"tZ�f��2�����.����>\P��܏�[�s6x���2_��ͥ/y?}C$Y�3�]M�R�ƙ�����b]�x[���98����`r�*g'{I1�xÆ��!#���G*cETj�H�s�X��^{�ޭou��x�3�dd��:F���Evm��4����������*k��X_>t)��ASW������k��~����\ffe��\�>mOCM���-hZ���B��j�����#��4��RW�03S�q�F�<zT����@�L` �}o�_ j�:�k˂��SIn�g$�>��^�BK_����jU;!/s0���wL��.Qʱ#�o�m�h�#�p���S�������Ƽs�_�ͳKs���xl�V�Q���...��o�#��6%��6��J'lg$��h��v�ŊnN14y�n���v\����K~�l���w
}��衵����߬�Ԑ�ƾ̜�^������b�J���M#T*��GGVƇ���橷pv)���(��3Қ��ٵR�t��R��/�u˺���ݽM�c����jj�em��ܹsQ;cG��^f�մ�܇�p����Co���(�29�4���vٱ�����#��n�LJ�s4�)�z�^�����U�Y���x�h���ԙ��޳Z��Կ?��`��p}������si�Ƒ��/A%����IkO~�-�<�B��j�:�LP�Œu܅	�C(���ޝ�!��.V�u8��٭d��7��s���Բ��4��J���vN��۷�޲���G����~Õ�D�~м�����=�?#�@\RRty��VG׃<�ssL�Ca��l���A{�_C�z+B�D���o���/'Q���wr��ּ*�{>.99fi)+לB��>  ���j���ȍuY��Q��`4K��\�/`d-a�Obbz��J�O*�1Q�Ū/0�l������x�����8�w֙���U~�T���*۫�X[+�{�g�����A*CBC�76�w����܀]�yt�r*BͶ8����{�2��T� ��ɴ���H���@����h�3�eJ�1�]ȡP�g��DRɩ�((-C/�E���%=�Y0a�{E�5;��x�Φj��3Ԯ�H��V�ٝ�F��F�qҰN�����?,�*p7������Z�^�&�sPc'�F�+��p��>'$�$g>���"\��Y���ݴ�������~Y�з8�ˠ-��^ύ���c,}}M�����<;@��~����+���q,e��<ڟ����� ]^+`z�Z�ԅ���g�G�i�<�$B �����\J�U
*7�Kt�d�I�t5�Y���g����]7OWݽ�(z#���4z�`�qQ˷|ٽ���|�Wq7"c��+grJ�l�G�X���T������<�+W���~?m�'�5z���� �#��\�y����w��R�c�V�桡��#��H�O�����S��bu��a"��ח��n�����W�2z^Hf��r�T��!Wt�7���$;�tQ@\�sQ˃���7d���^�@H�H��	#M������'S���e��ގ�_�F��섴v���[[ge�u�0�
��R`��&߼�5Y��_��:a������h�����O�V���R��j,�c4+��1`?>e_����1��ZӪ����9�������Z}0�؎��w�gG�X[[[zxȻT܏���n�Q��/BOWW�a�pCR_-	�������,s�[���P���qQ�#��3mh�W������o�3QSK����+� C_kK�]����s9��8p�Xe�F��hmu�-�܌8���/X��'Puzpy�B�e}�̤s�Y4���6,)W��MP����w}`	@okk����O �������<R>�uvI1r���M/��=8LʎꢧR�h��{	(ϰ*/�n#H�T�Ԏ;�x�����w�DE�ntȿ�LW�<ӫٶ�.�h��Н��_=��B��4���2��V#��՞n�;؞�1���T5B�\
m��Q�ɓ'���=}~V��t�5	�#��]��v')Ů��٤F,�trc%�%ҭ�~\1�tv>ەsY(==�▼^Bj����Uo�؇��?�6�A���"�5�H�Lb��)���:S@ڭR!7f*��h�2}t���y��'ǰ��V,��L�=#�t�� ���-=��4�F}�zn�ϳgϓ���ΏD?Y��(�N!ėC�(!��J���mo�U!��q�T�X�4Ə���Ug8Q�~���M;���� }�K��4��z�Y���ѩ�sD�H�B�����oD1���@�v��KyVS����hv�p��[�e��Nj6���j-��
(2�7d�r,yr�=��B���hԆ>�4풲��8��ړ`��.����.z O��n#��̬/�~�u�N���U�#3Mht����(H z�:0X ���B��-�^�$+ۮ��G���'~Ɉ�������L*�Gt�nI��P`O\0E��ys��}�k!!!��폷n�zJ)9�$��&M�����8�A��!�Gk[���п&��wo�[9w��~�]�y�MΡ[��=f�e���G�����G���_A���Uz&S��塊��z����S3��=\>��-T�s���G�o?�E�=}�4��bc1ף��h[�3��u6I�{��g���d��݇j��x��b�����o����츢�@�_u	������Y��e�(e/*IJ�Ex��CukgD|���0M���%:͉�]c,�#��mU(��gcc+x�R%��ԄGk�|nW��@`n�e�OԨ����ц����V��P���EF^;qQ@���d����lg|�`�#�sO�q��ot;�����b�O�޼����|�5UnM;>�qF�u{Jҟ���I��ƻ���/a�l������Av���hЙ��/G��D,�7)�rA?�@���1z�u_8Q����|�X�ڲ�a�)P��	Եn��5]��Ft��
��b ��HL3#+����#�^��	���c��Z�ǸD��%��_a?�m"�]�h͇VQOR�`��k�3�P�e�*]ũ�$�F�7
D����
ko]������Db�q��LM���F��H'�3S��1> G�9|���&��+��Y�?��_~���l�2z�Y��
���r|&h<����Ay!9��2��ʋ���#����
��ht���Lg�s�V�^�*:�bE�C�j��L DD�c_���,��s���9ϑ�0�ø��oi��G��4qDZ��I�gS7w���[ܾ�z�<q+;{.�Pۓ�a9�r��r����.J�,{���i�Њ@�B��	`�t��Fx��� ��Bd_��<wpV�c���N �O��;�t���D5��uv#S�6��(ѹv���|1L	�={d�z�0(���k�sjK�lq<;�>�D��j��A/d�  RE������D�x�6����ں�?���H��_��ǞB��܄0�(��ȁ���t�ltt� ��v\6^$Z[_x�`r[��_�����ėdyL�=o#� ��Qv��u���7�ޯ�����|(�X�ȉ)Y�&����_1�D��Ց%����'�y$V�5.1ѕPp̕}�d��("����y�)P<||&b5\[:���c̗���1��o�#�-��l^)�xxĉL�d��"N���R&��^���]��[}؎t�X��G��Է�`����H=e��n�/<�ָA�rRQZ��脠�F��� ���GC~�M�ڎ���`j��n��?�E �	��4>���_x�sB���?L��g�\O>7P�/*�
:�K���sn���0�Hol��*a�Nz���0�����	j����W��0��0}��
�rQd�j�P��� 3����V�]�QCm���m�����5�y� �����dp�
�)�ϟ?X�am���Tԁ�xb|����Ik�c��r�-t�t���R��ظm`��%�����C�)F�/������pF�_��� 7�㓩/=��~G4��4k	�Ig}%|t�X6�~�%A�=�;�s�����`�-/&	`�/���-ii����-n޺U���nc*d��uz�8w��kQ^�1uN.�Գu���-�p���d�77_�uo�tء�$H�L��Ҩ�y���3>������ƺ��P�騮j��Ww)S���X�p�o���p��E�P{{����i���C��*��=�SomⰮ�p S��=
��cZ�Mۇ�ŕ���0Py��p���-�|(<Ai�t�f�o����ur.�Ǹ��ݦw%�{$��K��ۮ������<��61{c�>'����oTTL����������b�w�&Q�i�h����/h�R�դM�s6��O���좗&���?O9-_i�by�@��4�H<�Ua���U������X����>��t&�g��6@��D�ĥu��,�c�J��9�K��]1���j��?�E��![}�[I�(��7�}J�m�w��P�����X�9y����S$�>���G�ߡ�A~[�"�)l��7l-k�u��� ��P��w�U������pp�Er��[�. �����\\\m+��Bt��F�ز>�����G^_���OV�_�������0x�@�?�Z�֧ǭ�r�Ŋ�i�tvI5��s݊�T�%0p����vyujzm�-B����L�ׂ�j �er����#@x��~��.j�@(��^���������g���vg��w�WM�A�}#����v/e3+�1�Z����wR*��
7ޖ��zz�@�x�nG��Ok'k�lA-B����M��>q������VC�����~B��L
7=~Պ(}��J�*�!1Ҋ�X\Ӣb������bX@��2~u}y�8�|�{ѹV�u���J����XG*��k��Fj�ZaT�������mċ�_�n!��/��%��zH��k�A�1fbh8N��=<��b�^��_
[ppp�yCX���\a&�(���׽�����$v���߮��k�+~�V���K��Y����XZA� �?`���Z�5�s�������wɊ����]��������{�õ��Q5>3}`�.%W��x�!���ah��ŧ��\T{�*�}���$�%^�0љ��K�2pŐ��<3N,��O�c�s��'�g���S-TN��肬�ᕠ�w4��� |���M,O����)�Gl�*ޮWbR��m��Q'���0����W6���^g��P�A�ر�sjk������Q_��Ovt?�ʣ���O��F����q[5��V�5wC�!��%��Zj��ړ��n��a�0����"��	ﾲ�2�z!<.V��qQ큚��yi^Ŋ���Q~5n<`�0h�����L
e���-u�����s[Cö�C�g]���(��"'�nˍj�i8oed�$m8f�j�K��@��>�Vy^��qdE���8>� A�@X��In�`W�ĉ�9��ų��A������.#A#p�}۶o�90�_��Ý��({F�0�9�R�t�'~Gw�W��C6�����AIi �yD��]���"�.�̶I�K	���[�������l��݃�XV�Rv+��&^M��3K|�p�V`���t�����8��h"�~b_PF�o�k׾ж�ܰ*�$�`�{�+D]YRv�K;��n���2�	�����(A�A+noG�pОm�L���G1�c������6颫$7R
w�������Z��=��2�"E���bԉ�73H��wڞ�G�@?f�=�yAs��?n�k�!�>���h�ހ�X�8����max��kr]ϲH��B;��%wG����l�&4�������%��}i��=�A�+�4QDih��-�1Xf�0��~0æ��)lR��;~�x�F,'H;���y���X1Z��ʅ9Wd������m����ce��un�^��i3�c��>�&��E��{��°����b�3N�<}������1>�k�Z`��\�]�^:[ƾ��%J=��ú�R�N2��}ى `t5�"�l�n z�Oa�xm"i�M>zs�c�	�:�1��C�)�o!�.�[�p*Wg�L�L����rs��~3HZ��my���]->>=���0{
ɋ�����<YɸP�'�}@^����U�jC^�y�r��P �����wf5��9߇+
�K,� �K�l[5�)?M�PĻ�٥��+��y���	lа9����2��9��F8���SfT��aO�o��0����M��"��E7�&R�+� �s��ǹ�1�Te�wnt�Ӈ�HF#��o�;�Hq
`�R���|����̉�s]&��g��T�t�j-�2����d�I����:R8L'zJS�B��q�#^e/���DgN}:�R%I�:�۟�{��c��?
I'�ʦ�3o3&��o1�o�u��sͼ���2��m��t�s/az+������}͹� �ii衙ϼ�e����/�*�x�:8Z˯nNB��U>dd��j��՟G�ج��n�x$%�K�&~6kg���_� �uݏ�����lEP�7�\��N� 4�ҙA�"
	���6�3q\w�m�=!�qκ4L��f�ƚ�s�W�a�h�@��T���f��v�4��n)�;ww���YI��)�|�����ҭ�֛_ �Oc�Q]�n&3�տU>+,��3n�	ޡ��B�k���T1Y�	�W�pG睵j�� ޥ�9}�Ѽ<<q� ��{��W���8`�An���@v�6�\��i�c�z'�.J[��fX��	H�A|o��Z��y��s�eԋU}��E%>��DbU���D����[�#H!�S5;�>���|���c�`��Ũ���D6�1s+����Wȭ� ����E��q�:��r�u{�^\Q�HgMy����󝬰�v�.$Ӟ��"x���%57����g6˝�<���Xa�*
7:�qfo�7�%�?o<,�����zf���I��},������^vY9V��	�(|ͭ��"JPE|�!Ӏyl�2���gC�S��]��T�n �����R��Q��S��nHd.Wx7�gʴ����릔�����!K�u�T���i�ܯ�X9L�@v"��V��K5,mЌQ"��1�x&�%s����wJ�n$(�
/TUn��PhGv�Q��OwD��?���#2д�h-Ɗ��t	�a�N�����_�hk��\>�Т	0{����g\��(!>�WD���@a�j�֕����c=e0Pb���3n���a��7���D��E��Q���|l�J��Ġ��u5���L*~�:�8��~�����3�Q^WO������5�@D~u���yp��Ci�۠Bt���Z��{�0ۆ֧l���Gz�~%����i�� 8H��H�#��~�^|�z����@��J�dk-��k�����)F�M�C�4�}%7��+���L~@�
�w+���$��{�	�~��b-G.hm/@�Y�����;>�k�i��nA,'%-�K(L~���S�j;�4��.���!xf�O��3.����C܈�����K�ԪydV��tݪ]��E��� nT���	6�T�Ǯ���St.x|����k����ۄYr��r���Z�x�O�KK;����Z�=U��!��>o�5��B ����69�&F}i�d0_��VM�pA\?��M�)�xORC�b���:4�dt�A�;�q�(�Lg���G��j�u}���
���5���9%Co�ْ'9fQ=`\��ߑ貕�Bx�4���>V��X�^
����xW� ;$f���'�T�k@:zw�$�����w���n����2��/�QJ��0�`�lШ_��K3�ɕ^�����KS?�L^2Q���:�i/��O�	nz'~��#������g��+�IX+S�`���/��},g�Y�����_a��F�6���]o�T0��c?�L«�z�8��zh��gne���7V��*�遜�M�Q�yc�5�'jo��6�)S<H�fD������_c��4�=�-6l4/^�R�s͍Yr�6�:���T��O���ؕ~E���H�6��N��8g^���T^�յ�z�13}�����1�A�N����p�Z�[���q�w���"6�̮����L^��Κ�<�`A2Ȉ��� �K���d�;drD?�Zz٩r�x^R����B���.']
)�������2��'&��~��Yg]@$��Uwd��n�03n��v􉶓9�W��1�����#Ji�]]]{v�9��W���7O9�L-�̪A�V�EX�\�;�:���_���lgg����MF{�0>o�Kωu�R�h��ұ��;X���СC~��8�:�}5r����s���6�O`fS�N..�W
�cX�5 XrL#�����x��XN���p~�U5g�<#*�W�ֵ�?���Z��].���P��P�������3k-vXQ�:�w0KVFf �i�].U���<�`�9,��}��կ�Æ��oq�,�V��Rҟ̏�Tę�1��{�n�:��y/�7�&^��t�������.��2US��X ���.`�ծ,���+@;1G;i�͑hu�ʂ�PԈ�o͐Gɮ���v���$�M�-��>@���4��@�<P�G?9�yk�)B�^��$�;���{3���[RR����a{{��6j� ��_��6n��5�+�-9N]���&����%O�l��J27��od��ӧ��HZ�r?��	l��m>9s�g���e!�I/�#N�{�m����̺�@X�Dk��7o����a '������=�����Q(	�RD�y�ͺ>Wr3����<jq$9�n����SR"2a�Iz���3�_v-�`'U_��o�ju�K��he']2�^����γVb����N�ioI��&��\�o�:�_Q-K���5�r{aҏ�9�5�v�ơ55��3�Y�V7	���3���ۚ���y�@P����|3��
�ؚ�Ȉ;���i7V�����\ju\���]�r���m��!�9��=�$m���K����ls�f��'b�(Yy~olM"&����E��.YKٚgIJ>�7{��dq�x#/�������}���F#�����m�zc�ן���<���A����|�ԍ�F�k|^�p�om�V��Y��Ɔ>���!L�JNd�u`t4Su3��*���qz�� D��y�j������8l�������{э��0sT�K�D[>`4Z��m�Sئ���K�b�f�L�����K�E�����9N��&�c�s��(�^���2����$g��P�4��H�kV���G�NaI�,����/~+��U}�<��+��µE 1<c���ߝ~A��[p$ٸT�8p0~ZC��ew�V)�FB��o��t�  ^���A�.d�S_��8�Ҝ���-�����vϟV�+Dtl����XI�Z�Q�<��q��҅��ݎ�'��H#�& "}�=�9͎��y����j����@�e��@q[>�b�{Ĳ(�
������6�K����H�?.������M xB��q�ѓ"#1���T})����t\U4srsŻ���u2@��
��v���nf�jr$]*�|��oڹ��o+6JWbo��G��xV�Nk�� n�H�%����5��V�S�MNճ>y�D�)0���ř �{��]\\|M�m�@_;tSV��9�#���|�W��r�Q��^=��^}�2cԔZ�_��MP/}�d�g�넔fh��I�8:�_��3���/9n�Sui�n������F��O���^�*)qD�Y�D������㕌�R26���$g'��H���'�#�~}z~��������e򿈈��JKJ|��u�H�u�~u^���H���6\02��)����T��n�[�!$2�8��겚�k�
�=��7�.[��Ġ�h���h�A�r�e��=�x���I�/B�9��%=�[�wMїsvǍ��z����C�;8W&�@9�Q�ji�������~�(}%��g�k�P2�pƝ�����n�a�5.����ʂ��YD��Z�_��,�@�{1�Y����K~Р�:��Fo��)��':�&�g����)������u%n�_"Z����t�GS�'*�9�0�4o�-��5(��ϋ��Tz�͈��{���J�(�Yj�.�$Ž�_��4�4kd��&0R�pj���1z��Qa�����`,�q)J߻)6v̙���j��H�����&��S�X�T���ߏ��XԄ��[]ȹ?�,�����;����s��C��$5�ǩ{���^K�������/��ء$*#�)-++ہ�K�2�@� ��Q�!7��xV>���-$Q*%�-R5;�C)Y��zbae0
�}�`)��ۯ�
�Ǐ�2��{����r���Lė���X}��oAB	J���9��[�Xc=3�b��\C�<֊lJɪ��DkV���U���-�+F�)����yx����� ��	�KO����,_y�'DPz�B�'�ka�9(9wDaҶ��ާs�`�5����h`��Hp�zK�vy�:z��'�B���_fI��1BH_�~S�s#�A,�����*_-����}ɹVܥذ�}��g�n;����b.�<I�^f;���+�z�CTSH�{S����ߴ(�,������C�3l�M��U0Ӣ8�XU���2��%n�;�ʱ�����  {�"��}]�2c8�o�^�֯"�wu>_<�b��j��7��(�|���4<�ф%a�sw��J�Y�b����Q�&�KjE�Z���j��봜�Ɯ���V��B偘��7����ʮl%V(�<<S�����fF�KVv���V�T�Ұ��[)3#���+-�>[�ib�^Y��&�LI�`x������eRyAA��?y1+}N{)�^��:r8D�[rgg�f�>;�qb@ro���dRZ��yx��ʟUC(��+�̤)Ig�=����ة�k����qXM�8ݎ9��r�d��!�b��}B.t���:�t��{�[��}T/����'���!�q`�eCT��޽{�m�sl����K�<�a=Yǽ�����\&]�f���\�#_�C.�n9�Wb�|��K��@�/P]O%�D]�|��T��+��𜝏�ȻͦT^!&sC��w�:��r&�����L;^+���Q�㏼D�af�(B:�%�4�|�5�W~L��2���~|�<����<L.����Kt�kӨ������@�;�N3�x�a��VG�r�ZWW�aZ�Bl�S��r,?�J�і�� ߝ������W[!�Q���2A�@E����v��C� ���nK����)��+��UA�-Q"�hʟ��i9�j<?��P��r�c~&��)X�>�mb�+y1-�uy�G�2���?�N~'���e	�yG�,i`- (g(����FL�v���ըC-^bFV���C�}�Qa�|�^�!TA37d�i���]�*�;�x��5��Kr>��st�ԫ$N�sIMʴ�Ӭ��u��ϭ�6X�s�u���8�����(�g��c<+��8��9:�z�m�.�kb'm�صp�t���Ȉ�n�D;�׷O�F�=��Zk񲡻�֚*P'+i���Ǘ�+&K����j.:Լ�R��Y��f�Fϔ���F���r|kW����C�(}_tb�n�^��� ��*�V�Xi�u��)��@�q�M��O�m�����P�C?���q�� *�����)�� k�;n��p��!�*���VҐ�FzR=̪��`�2����f��7z����Ml�5�i(�6社�s@G"��W淾�`���ذ/�ᚗ�^"F{�O����P�� 2��tM'�J9Č��vs#0�{�q�<�k��i|?v	��PMO�?�Zp��&�Ss��.�ڗ��j\�a#!�~�ᆫM��Ǡ'{�� `�`��Bj�����>R��$'� 6<z��hW}}}�[$T�ؿ�%���.\�*T����J��]ϗ/���eW��j�E3^���]J�`o|YV�x3�IKK�r�#��֯��3�uW�̖�Z�A�n@$	�IhI{�^�tV�R�y�����ݡk."#�(隽%J�[�l{�އ�\�4^�ٞ�����|�Fn�����$'���0b��ŧn|_��T�
W}׿B���N��7��Llj���Іt�A-VB��}ԠO_J��*�3=���.kU�����[��yՌ;u�p]d4>_�V��5��`O�v� `Cqׂ%toÖG�s:��I��@��
�w��ڧǽ����H'f�����'r�;�;�4J�7e4�)��yR^��?タymn��'���p/��U�2rOU�9냩��J���K�"gZ�WYQ�-�6�W�}|��Į0R ��f̴q&wCR����ѣ7�!��h(}��+����Ul4��{��E? `M압�Q������ڢ�.�������'����i���L~��lx$p� VUl�Q{��P1\͈J�+�pW��o� *i��/ۃ�l�>���.q�X�Z�TF:��^�ȼGe���<w���q���ku'��z���]B��M�ʡ%�\������8�kyz���3�D)`H����6@����23���.cͅ��vX+��i� '�qw�L���!��z�!]s�BS%LO�&�!�a��v�}��̊��ZN�k׾V�׭^��ϣ��M�
��h��9��?�z�ҋ�ڭϭ����nGb���~�d�Jh�0I�rD-�~&X��MoWVF�WFT]G��$�SOSS�s�"L�a����9�G�� h�#v���m,��:���$�!�9/^��?�N��j�Ǡ���]i��'6����q�h8YG?5 _m�¸��>�_YD�s�qh��|�=]Ϩ��!�Y�b!�����{��88L�ϐ`�.k@{d� [�ێ��޽��\p���gDFnC��{�v��$}��KzW�gX@b��<ƒ�އ�싻�����u�:\�H��KƾK��T|:�BN@���:��y�t-�1�\,�����`	Yd+��=ܓn�H�U7��1�����p���<Z�lF5m�^�k�D�̑��Gd4Vi@�F�}_���0skX�5�%?�g+:��DV��'�J� �!��f��Z�r���Nϴq��7���X@�z.C#0�̏��H�����E�r�91I~:�[��?z��x�v��:�
Up�)Y����`r^+Z�w���O�s�7����S�f�N����)�ރ<�)�%#j��h�������AC�ЇҪ\�'ˁ�H���߁��`�O�1��W����C��%N·f��UzP�ǿ@��P�墓�{_��\o�?Wp;hVI�����Hn�/�T/))AG:I1�_�nU�M���B5ڠ�hL(�]'>�'wu��1�A���^�0���u�!o�8��S�ndd�v��	�]�������-5o9�&S.Hvt��u�(��t_:��vh�H�K�9=��۠
W;�����,>9��n~q��jm/R;�&tU��Y{e���Zs߻�Y�yu�q��VUb&�9r�"�h=�k���+A��.W��B.���"p�j}�}�_�i�>�8p��sjI3�.h�o��te>�?/��N'8!�ov�f����ʸc�9u�֞����6�\�[��?�]�Dñwa��ݚ�yϫX�S���e��7op{���w������r��Q���7oޜ&\�mv��Ә?j#�B�_-�{_>'�*"�����������Tty�DI�(�x��ɚ aM񋐌���>��ϸ���\;e�Y�1#�/l�:S�5F;����^X^H$����?3�#���s}�P2:�J*��ζ��6�D��ڳ��&#j�垿W0�Y�����.!�����~ן����v<cd�K[D�)P���v(���c���,����(v�'�Z��
�Y=D��c?��ͺ=b�Β.Գn�	6�{H�BK�Pd�h9� m�5Y4ck!/vp"5�L�Z�p�#	�@�nAГ.󔎟YD�ZIE�����K'|;�#���f:B�wF���z��쬄f� ����B�D���1��zM�vL�6g0��r[�����0���	,%�6�:��+���~�^'����ַ��y�Ol���w�"������V�v3�D����S'�����999���g�mb�z}tb����c%+���"_��%�e����-�yé-�\A���j
~y@BV<+e?K�:�>��]16�݋_މ��ҏ���UX��m�iZ@[��`���%���%%�GC�A��N�j����]<�[�L�.��~�׀P:��F�x_S�֢#�P��$�F����I7�[؉���kRn��T ]K��B�0��)��Ϣ_��~�W�&#+[}#�x���W7����ܜ�㇡ [ ?ֶ9��%�ݷ��[ODT��Je�H������7á�s�%V����E��K=�j*�g�5	ߜ
��)�����S9��񥠷��1|��p�����En��(����l	�硟�F��o�O�N��~7}�&yA@�3^�����4�郞P��p��Y9�GzzP���+.~���}����nk�W_�N��?B��;���߂�j>G�W�Cy�̟�_���d-uX1��`��{\��c�Ⱥ?/��g!�|G:	�it����x�jq':��twÜ�L
k=oߞ. ����R��m=Z6�`w W8$��믥�(?��$��?���9Pp���H�����Ë?�$�+�nz�4o'����6hl[��itRˉV��0��̏�ƐY>���
-�N��+�d ++�Ld�s9}�tr����g��j?~�H�ƅ@z>g�v��u7V��(R��3ɲ��Yi$)L/��E�eu���B��'7�J���ݾ
0�]�k,$)O���8�v>�f�w��6a*2�f��t]���V"�	3�j������WǍU'Z�<�]���w�c��ٮ��5dP����P���f�z#�]���y������%�0�n�7b�_��+��U�6*:�/��i�f���O�A�������"\�Z�ZI6]�������f��~E
9/����(��+n�*w� �.Xh�DA�w0�{���������k�BQ����[���w�.޳{+���j��<Ǟ�W;t���)��]�#���	�X������W�It����`��YOC�(���#TI�?��;������3*���q��b$�`D�
R,�:D%*��P�m�Q z���Hs�л�J���;�����?�g09��}�^{�s��y����0��R��.���C�:F���ky,���������|ӫ�7l���,�����j#���8��������}J`!� ��n�$�j���״2)�d��-������6����B(��^\��ҵ&(��Tjj�M�;� �4 £ҕ�c���>�{��F;��(P�]�����VƦ�1�Abo�>�R7���cUzi�b������9�)DB�lQ_��H%�F��vU;�؅?��c�ޑid5|�ԑ��^ �U��DD��9G���UxJ=K�LG�`����x3W�L]/��$.]1��	õY��\��'��#F0�W�2[����p7��ύ~�*��K,U2}�����f��X�2���=Dz@&��<��~u�+X�/�X��í�?ݏi�K`��B�NrC?�@����"lM��o#����HD��#�������^���u}�k�\�����U,������qo
�ajS�𠻰���Ti$�"�f<�a�:��@e:v2|�3�;Us��~MSǪP6��4|�)/��A+sC�r��ז.X~ìO��y�s��������:X�Gw�ݸ�gJ��߲�v�A�!���]\$X�ښL���^\��������V�ӳW�nmc�]G�dcx�V��qǐt����"��r�)�{����~���*��5��D���]E�WݣY�n!���Q�W-�M������W��pa0�SS���;`zƟ��2�o��ߑV��W�z�a���T�4��Y�T�<�#e#'��*w���"�տ��0,�������M�>�)�ǋi�88�ﮘX����M��M�R �"m!=B�B鯖HJJ��vbo�������3�F\9]�1�뵫�M��(b���/� �7����w
< d�.;�=n�C=O"�-0�O�>}��ԩ�=d�-˔V(T�=(�"\s��Ks���Ay155ݷ�$���gμr[��ҥIKό ���c�u)))V|��b��S@���~�$�Y�Q	A�zf�ŵ�o���*Ў.�D/�?�8$*���,)E|�
�J�N�j�8��ޠ�"�%j�o����ɀ2�crL�����P��W��\	�>	�s��b(���F��u��n�惂����o�cg'���@������R�377Ov��ɪH���}}��N�XD��?MN�r���-�z�������i��Sc�^(	.�[��@��I^ЀUJ��h����O�� i�~�wr>h1	�%+���+����y%���ϑxԝ�����[�`:�DB9��+ 
�Z�Y
���gd|Ϝ��V�<�нQ�Bi��ڃ��7���y+��.M����*����J��@7�>c�&�[{Ztq��?u��������Ҳ��vHW6����廒LW7w%e����R��n�tO�����`��C`�9.Ns?��H�l�"i��>�N����)C+�O����'��p�e��_��*GRx3�LPV�}��Ý0�1����
�s��� �����dg��ݩ���^�Cȯ���6l�I�;c�+��lI���*a=�N����J&&���]���~�p��!�z|k۝�c̕CX�L�^�U�g���ݲ
���xiD��Y1Z�330S]X�2��Q��C 9����lI��$#a%k *�c�)G��Pk���X%����=��=�$���T,@�.ɩ<A�c
���Yg�N'�|�u�i�r�#Rʀz>�17��y��n���!�qgT�ȄZ2�t7#q��{���qRx���-�/*?ӥʣ�	���9X�6qRH��tP�;�0�<h7n/����-�
�G���	'�	9�p�P��Jj�W>�xz=W.�tED,H��Y�q�b��}����b�P�i�A4��hP��)T �p�����b5.~[d��'*ߙ�� �^�-uv1\��A8��W�5o�ׂ���m��w�K>��z�ξ��*q� �mu+�����?�-N+�����t"5��=�/��իI��#\\]e��O-#s[�G���[�#rW�}T����{fN9�<���A�Ǧ�A��CQ3�֯�9Ԕ��k}6?feo/H���p�W�_�Fqt�fD��2�mԥ-MP 22k��A��6���"+�U��E��Q~������-��+SYiu�4���p�`:.�h(G�P:�	�LA�,��K��}�Ľ�����~w#���"MtoP.�ך�A���e�������swR�r�&VcS�ͅ��D��o�J��UP+a�,�X��2(���oܯ
�an��;=�h�(��t�)�g����H�d�SיA.�G��B���Y}dsp�3���%y�Pڃ�1ꀥ�� �p��!ٷ�K�� ��``�Q�bf=�2Ҕx���=�s1���T�.�@Մ2�%�,�x�QX�B�~	?z�J\�k_<Ճ[��(��[L�[��F�aѭsHˈ�sP\5��ǜz�p21ȡ��9A�b��t0w�ӳ�C�Df�E_g��c��k�!��E�E�KVR(��#sT��qJ�&���؈�׷��ݭV`e΀�;���N��"�yx���_��\q���gE�B����RЮS���@Xk!����P��;��+?ruq	�Qq��(�Mp��
3�+6j�#�(L��y��́��Nl*�^�?ѿ QΗ�M�v'�Հ��;/b˄?]��Ugg�]�N-<��z`~�԰P#�0��6�:_�)�Q�~�������PYJ��V��ҢV⤶H` y�[L�4�Gb|V�튟�Ӆn������Q�n禉����حx�9�L�s[�\dPQ�" 4JEK&rm!o��%<������-_?|��<տʠ�U��'�k��D�i��`�@qa��͟�i�œ�|M2V�P��/_�y�HF��������V&J�֚͛��MO|t;�#�D����#Em��+��]8��>pu�z����YD�Z�B���AF�q?ݒ�ϫ5�4��$��`rې�6ʲ�������]��E��p��l>��9uK!�Y���nNؾ�DDF.��\�(��t���1��Y��>J7�j*�`O�qxOq���2�S��sH�t#���Ur3X�;H� M�����
�!:o!��zᎺ(��	��'��׽��e�Ց���+A�?�,�YL!>��E��Q���[�f����XƁl=乸0?�!��["L����9��
nU ډ��a�/]�7Q����<��#B�ŝT��ݭ@�aK�/1v��sBQT*�B����q��lE?�F677w��_�o!�$m�bR��l�����q�Peb��~���G�Sp����l%.u]�L��xV/���2�{va���Bw&�9���-�\�H3�W�\������j��r��rBI���}�s�a��`�Iz��b �'���u��x�>Q���Ah=
����~�/OED��mp%��B�b����� �ٜ l�Y�d��+��zq�ዎ<��i�F���#�J�/eD�<��u0���2�'�!�@�^������c�ߑ������@��� D����Gc�q2�ᇴ�R��f���>4X����H�
�L����84�xҭz5��/$Ǣ7{�Om?��7r���;���8��w�D�{<��a�����	��W!���G+3��H���wK��RV�1I�ktD�97b�b@s�]_�G���Q����Ã̺��j�F�P��BZE�7*W=�B�Ǭ)N�?@���}��?�)�MΝ�Y�J���8R#^@L~V�v��-��B@�I`�" z]X���m䠯���ᑴ-v~�i'qZ�K�a̡6~'�
��)u�3থ�H0a���������ƻ����N��ܿY�=����`SŲ`�6�`Sf�$i�@�L��{;c�̙ˎl���{�9+����?S4��]jb�y�:�ٯLԞ/���F�+�������b̽��Z�\��v��}��ǐUiK�A0l�/�����b�޺�#� <��HI�D�'��� ��@#��oذ!��O|BD�.��X��!��ax���ҫe�k��NT�ĳ�-�k����TD�2~��b�45�C'84��H�j�koޟ�M�ɾ���Q3��R��k��P�
�;w��"y��K� �y3�f8.}m?Z?���R:8t�)�b����ԩ���;帀WpS$4p@����Q$�zH�D�HPg���lGՔ���L�Up�9��߼��)o�53[Yh�9p����#*�þ��x�*n��x�������[A����Zg2��F�[��Z�WX�Ȁ�;N�LTS����S������n�'.fgAʩ�/��B����Fr���ғY�c�O��\�~����@��V��@�5Z�P_lf_f������"��>�s4�����,��b��\/��讞��7��/3RP8xA��'��͗�o���.E�ϻU���H�ə��[�j�6��*Q�įAߟm�u�*]>H|�L+��j[��3\z��z_�u)
���	|�o�mb�s��XM�D�W�E �o�+kL�EjQ�� �lg��DB�8�ĥɍ���W��[�8������w�|�<H����-A��/ޟ����f��}�^�j�S)�Y(Ҟ,����I��2����:���:�#���<���4l{
�Z6g�ե��F��4���9Ků��S�Ʋ�7�y�*{/xYz3%���d�v�\ڶ'�.�%��L���>�W�?�o���"���q��('�R��R����:i�Ny�ˑ�X�JH�\y�~	�ҔC����,�o~O�͛�e��d*\�#E;w�:��C���l�z�0�E��Yr��G?���s/�����ٗ��J&��Vimi�Nw*ؚ'`�I�q�z��fNyC�W�|��k�Xzۀ.0ǚ��D:t�P[�W�Vi�E���̝W��)B���r��tK΁8��
��Q#��>��N$��2;?����g�>�wV�Hv~$y�B��]sL�5+W��bs
��e�,����d~���y��n�}��9`G�O�����Qv�dXeE8C����9Yخ#C9���+�B{k���ve�4����H���:W�ƖmR��v"D��|� ��N~T�|VW���>����k<���" ڟual��`���K���Io~���_AE�Jy���&v(N�6��}� �nla��g!�9��<΢�jK���65���W��B�9��.7L�`N���xБ����f�z�4I�V=$͵�d�nٲe0�� V��8Ln��.�Q�x!����@v� -'�j�^^I��HM�Ӭυ�A�X��V�@�差_�fy�}��	�����4���B<
���Y�6��V�©��퐋���"f����Iĳ�ɝRi�ă�����r+�:�BCj�z� ������ۙ��:]�.�v��k�e߹
�G��=x�Ţ����������hH�^�r���NYM�)P��jjj�n0���06ȁ5�_pdO	V;~������k�l0�&C�T+�wD���Ź�s% ��3�M��Y��ѕX��q��q<k,M����S#����W<�H��
���899�:���V���=U��-F4�a�Y{�SJ�ɰ��d�(��т��10a�H�G C�����t�����y#��"Iu��vJ��יu�%~�R�>�������1�G����-�⣋��>��-��H���oϓdג�@=I�	_�t���c����dW�'�P�-f0��эFFF�o_Y[�	�{��	��W����o�&�Fn�:J~k���H3���� &&����R������z|��OTTT�����x��iJ�o�ߪ<������q�9'��w�5L��=��^�4ʣ
H�-B����� ��(x�l�Pd�*-Z��'�8 �r��k�q{�����ǂ�u�=m������lF-�ug�?���c�P���{�!�s�ls������΅�~F�%rKxIz��2���6Ah��ܽ{7�h\@I{+j��y���(L^Ԉ�����=�9�!Y�"��)(k�OTtڮ�^e�)�j(�<��j��g�� �(�>�Xg��������ϯ���y�Ef'�a��=UB#6�nejC�z7�xw5�U�Ԓ[Ԓ�\³_!xC�F �U�sWQK�c�''8�w��� z,��ݻz�p�GORQ"�΀��~�MO�
�ȸͪb���7�GH!I������i��H��˅_y�-oy��ŋ��'�}��(�Y}�����+p� �%��&��/���"҈R��ACVFƧ�0�k8_.���ԝx�@س��@��SVV�-.����p�z����%���9F�ra~�H���)�J�/�U�ǏȖ$N�����SE��mXG��:�sZ����>on���Qp����T� �`�o�cb4)�|�f5Qw8T,�3�N������7W53;{��VVtK��@����Ç�]'[���l:�$�E~��`��~�t�20~2��� dIz�Y��*�w@�Uz%rXU,�皮^�:���aD��8�ڔL�U�q�ι��**+@�?�D��-Y�e$����ŝ��X�ɭ�C@�� B����;a0����c��¢/T�Z���{��{(Q�8<�����>����S�u�n-�[��;|xD��L��m��960h������f}��Z]6�s�H�ZZj)��~!o~6k?J�_`�oB袓y�^?:kTI�������&$$�F
qe�Ls�^]�(���R
�˼��p��;lJ�F�ts�%���탨v�ƞL#�Pu@���Sq)@�u�QXױ���+{	ն
�&�;�gp����JX�d��jn�8��W�\er���C��gv �KG\ߣ9R����fef�g@~f֍��ui��|�(�q�R?uE�p������P�+I� G���e��?�u�+^�vS�Z3�f��EGvk��J3ss�u�W6s�?�I��a�]A��9�D<���{�QX�n���_�par��<a�S���؈�
J�Y6"ۺ]Լ�Z�b(HzU��{4WX�N�j	w����b���$s���1	���̤�Rc������>��kI���¿��N�i-7����jr"�]SOoo���c�Ќ��4��A.D>�2��+k�2Q�����W��W\]��^l�pΔ�j���m�B�*�H�r[|s>db":5�y5p�q�)l�H6F�w�&������?K,������vbJ[Z�Y���k/�/A7�r��7�ڜ�����H�����ȝ��34��s��d��Yii���N���V��<��迁��v�'��?t�8�#!�3�M�J\􃃅��5��wC�[[a:Lօ4R���]�v�v���fسP��k��L��A�Uk�Xx�I��D��ߑQcH�
<e�4��i�N!�z���~<�c�#lX�b�L'�����{���x���J���ѳ��+�S-�d+�xeK��,2�9��N��6o�s�
����_+�p��������4R�[���ڷg��95{f��\r��N
�<\��?z(ܶ={���z/����q��azO�n�h]V���6�P777�?5���GVn�̔�~x�ɨ��x�[#���B��Ke`��wp�����C)�%��Z#����N %�3��~m�ǉ^��)��eo���4�^zr��=e|��5��|�̠�FJ,�]�"�C5���}�5�5K0b��)6^� ��<��;(��7��ٙQ]����jei����m�sPw)K��É�7����QS�l�'q"���xfI5M���������o�)�E�`XeX�0H)�~�шς��;e�e(�f�f��=j�Z��o �wv)*j+��,�yL�v2��u�=j��4
C��7�*CҎ���U����w=OJ�;�3�GCB
g���}�˪i���ϵ��4��ݓ�	��U�}�|M�B�K�"��I�A���,1n&��KSs�_� �D��so�M@�CUcd��ۣ��Z�Kh���,Z�Y�`ӹ/�q
5�D^���IYf�W�VU�ă���r�w%%%bԒK��3����a@�h�Z7/4�?dn���4���/�^�-Z�8�i+��~aFU��/Q������s�1�M �����pH5��)	'%%%14l�. �/tB��~ # �W"�P.(�(-�ZWo�%Z|��a�cPѢ�#ۭ0�������ΟE���[%D�{�RtvJ���-B{��}�����s&N�lR��f���Vj#�	@�
�fJt�_��^b�������f����YR���5t�Dx��RT(_Sab0͆"�G)Z),�!܌c�?=[o�[x^�u���9G����.�����ɇ�_�\�3����2��Ȩ��#��v*��h�0켬�c�5����i>��2r���������O~<ofW���}�{���;w�.y�!/ό�p�����>Q8Fr���x�|$\�|S��qJα� �� ;�U뭕��Y���Jy�_��Z&��[?ۀ��!man�o�m��`���tFx�c���l1L��_'�O|�	��iד�&�}pҗ@�*��@���KA�xG��ߔ4r(yG�^�U�tyB�5.7Vkfe�>�oE-��������"<}�c��&�Xli�낧7�[���2)�@���Osdg�}e�ы���4`)EZ��o����8?Yt�̙3&�T��1�vM�g�X��5[�ju�zw�(�xFE�%��Ve@9b����z�/�0��5�4WOF>����ҁE�%�VV51;O�
��B�޺�ufVP�3^�L�7���_��whRL��V�jx>E�EX�#Ti)�*��;��N�LKm�T�p>$�%��C<++ַ�>�SL��P�b>����گ\��!�.�[�*�k�+���Cp���dKMɰV̸�hW����
o*��ܙS��!����ВZ�X��7?nK�G�Lbxl����F�����ʬ|gf�(A&w��������'��h��=�[z��<��)|��ķ39o0�:�wԍ��/�V�ރ��-ya�{��9��+k�}����F"!#��̬<�=K,l��3�+H'���Ƃ�2��ԅOh��u	#�{y+��I�s^d����p��
�z�>�!��������)�S�sG��>�#:_ݙ��=�n�@��S�O��.��w��.1�H}B���K���dwi�t�G=���R�=�2��ߣ�Y�:�%�I�rG��ϩ@�����n���
�?_��i����x�-^�沦��H{�����H��@����C!g�ܣU*���-���#FFE{�]��7����{@��.)t;`���+LB������-�WW
_�T$w@����/![�l)�&�|h�-�5����X���@ԋ���ڿd�׽�LI�I��$���>bae����a� ��w��2<|^c���/�"�oOe��6�y �-|�[�tch��S9s�?}biW�O-nPڭ��K�ܰ<T���EmE��A
p㊞���������=fS��\�5��͛�WVVN��z�(�+iDo;� �H:�$��^ā{������`V� ��`9�I6� a��:yN��K�jZ4��zlٲ�R��ij�cTԶxqDr�����7�.{���U���s�c�˨��sl 7.rw�S�x�:��8�O)<;n�<W�U����7z���(��Y*m�ӑ�f�F��i�&������\L��n��)�*�,�E�^�����&'�F`��_�::~�ĳ�,s�--AR�$��t6��� �X&��U��&���A�pHc��V<n�:tg�Lf�CF텀C*;�8�G��"��0��~M|�P	��v/�2{�9���G�S����)��}�;����NL�����΍���k���� ��9��ݷs�ab�y�
YVC����#���ꞟ�J�g�ey�
��y+t�g��h|/
���&����v�?�k999� ��X��V-g�͞��t�$�p�.BX=g���4R[-|E"�o�7�?���/�)7p����( ��4)g������� |@<��P���aNu�K���C!\�i�8���c��Ω_�N�XGj����߿';��J<R�eeY����y��hİ&��o�tD�E�@~�2��`Q���a+��<��1NNIY4��r#A���L��@9���Ņ{�Es}�J���9pOMm�x�$��$f)� o��U��dT����"������.Ϩ��}�D+�7�s��,�㩌����F m�SU�~��{�.��|��,��dl ��0�6J�1�B����O"��h�.�p
�,'!!a7���1�E���U��a1��㩙���D(9�ImCVp{�b�9��`��* ��U��!����۠��x)�-s8 �{<k�+��B��̢�9��ҫܞ踸��L|�g�tȯK�Q'���G���A�Y^'�����Mg������^���s���K4v�uh�>(��q�;?�{��P��.k B��L��*���~�u7�<C�}2ӹT��,Iz��ƨ��
�#�C
)���e���m�0O)�����5j�v9�LAV���9/=�mR��

*��_Ak�#�(�HIe,��*�(}�4�zʠ�!�a���%���d	��(>a������R�HX�SS���PRU�%̺"h�D�f���'�o�6�w�QƘ��0!�N�(O� �< �g虝:U�`�ߌ#{\���N�%�,�"��r/�@�R�h�`�|�{2�X��c,XS�t�s�-.DO�;�'s|I���R� tܣ�̂
 �~��N,�4� ���n<6Ч��
XCh��JRҊ����U#�rR����JBB�	�R����d��J/���������>9���O��**��Kn��g����h�~d���3����)!�	� ��f��T<�鐂"�mR`Z���o��EUYY��nI:L�����0Yqa�$����d.��j%q��Ϟ��T�fNX?E �@��9�Ü��[���d�W�iDR4$eE�.q�_0*�@α� �#S����A(,�Y`b,7���������W��=��	cc��(��(^n�w�N�,�d��R�Jͱro(hΙ��%r�S@3��\�R7��r<��!�I�Y̸�� ޓ&�ǣ����
9g'��ե[�IUx�;�h��tl�+z��|?�9T9���o������G2��QM�)�𰧳=J�	�A:}U�a�;�M��1|�K���Ӛk����! ��ng
ڇ���V�η���*t����}�R'xG�\ ,��Ϧc�H�^ ]f<�\+�`c�ԡ揢ʵ���]|0�+��k�����L���T�����z�q@�9f}�Ai����.s��(P�t���GЂ���
�)B�<Z.���L#���
�� ��Gm�)}@����g���C�B�� /��7v�oN&��#`�±3���x�5� dԤ���m��j���/R&��_<~p-E91��ehe}�F,��zR`O}Kۯ{��|�f�.�fzԞ4�o(��ʲ�����Rf��m�B��X�g�ղ���"�n5��|��Gd>�*����x�����Y��wk0�.Ő<.g��G���9�5DL.h|i�E'w%J���8�0�P��̶*��;F�����`�T��e�Nխ9���!uR����p{v�qʃ����F?(.:�b:�9�����Ox\�Sm�N��5��DR��^�{+E�<�)�ngx�H�����q��Cւ"b2�`�~m@v����` 'KK��ڧ�%�g'5r���Wlj+//|�����]�+a\i�/q���[QU���� ����.��8��y-���W''��~�^��w�<S�y�PGƕ[�/UE���O٫������z-���k���t�9��6��A|�I��-}���ؼ�� �x'+�X/������Wy���3���ٿ�	�KN���L��5���ݧ�cۈ����sf�%���#�W�f����*����jY��ޟ��6ĳ�ҥ�L��wk�B[Xs(t�u}ljI0�D{v@1�},&�.ށ��ؘ����b)&�A/XEYy�t��E��J�㧆f4�,K&�X3R)p�0ql�V6��nQxx6�l�{Q�"�7b���b	�`P���:�i�E��5�,|���Q��S��`��N&�g�aW�Л�(úXR8���s˸�e�*�z�X�p:ef������97�b[��fF�>����nQ�#�F�0z����G�B��ג���{�����@�تn��?>�τ�3 ���t
O��ܕh|�:[���	�a�ү�A#�����b>�� ���h��o�H�6Д5��i�D�C����篬S��>���%�
�s�����@b���������a�ٖ'P� ��$i$	�'k��⼖O�|a��/4�M��6��)��s/.�Xb�Lb�^I��r���A( �����hZ��w���;+7����Eu����V�4)y,Ϸ���?ȉ
6n���EN�Y�#$h�#�S�j�hB|��l�@s�ۻ��%ؽ-y�:���̩���(iikq'h@-Jt��тd�婫�ьAI%ef�LdL�����s�K��g����!o��3� �H��Z�>NG��K�r�}����u$�� ���K�"���x�'�zq�����das��uv�����, lL�ʫ��6I���9���ʝ�M��q����K?@�o����-�G��ts[L��I�ʥ�tFȧ�^1�"�5��Dfj4�.袸�dp_N}��I�ۣ�������sOI@6@15?�[R����'3��q�� �L~���*XU|�)�y�ש+ĥ�.s_��:�h��S�L4UՅ�=�ڵ{w�9�}���	ME��j A��c�ς��r4oSG-�ǧll�j+��r���(El`м	ŰWDN��_�~6
e�棸�B�Α*�S� ��`q���T$O�#	���d�&�J��kn�Gǽ���Ʀ�����z��\�hS=
���t3��;: W� ,�=�#خ��:H�������dţ/��r�{M��x+N@�XVS�{\D�	V��=�����W �U"/��i����P��0��5�$@tk�~���]�S��L|�W����C��~H����$�$���tzP�b�Y_��8��s0��x)|2T��/"�?���Z)[�"T/;�7T�[R��� ���ڊ�����I�0�{B"�%
� ���/�$-
+P�i��I�U!�V��[�v_�n�����E�4b���0^>�F���Y4M�K/kmՈ&}�x�F��fj�l �4��0�PT�]�3�e�O0�n��Z��^�k������#b�_��,��Sk��k���񙲳ˮ=w��HmR��h?�ܿ��j��9��,��X�&�kM��5�Uđ?466挴��]�ϔ�4ǐ�t��ݩsK$��W%PC-A����?�t�ډ(0�M �t�Xt@��ࢲ�e��w�Lr��ӫ
w�� 5�}�x���%�y�,)Z��q_=`jx�M<|����h#�2	�Gd� h�ªfu���KyV$�k"uS�mό���~���!���ٸ)�t�$�����]�R{�\(�9�g7XӘT���0E��%��w#��"u~�]�NԘ��/�!5y�+=��Y�B��=��>����p�wV.M<��q�Ƈ๹6��?��j�^G�k/����<�!����g|]X�}(����X�fX�qZn;����h�_��	JTp:������S��
�����a-ԇ�[�$�ǳ��ڂ�@ޣY�=�G^pT���,���32�onn�NC�pä��1����[�(�@\փ�ȼ�A~r��	�`l��!�M�b�L�C�̢�_%|�A�;��c!��oLTO܃Q��%��s؈�Vv����PKHH�c��V�);ҥ����f��o�m���$�m�}�&��#i�{ >P��c֓��	�A.\7���5�My���ߢ�E�fɣ݈Vbx�S Z3��T��܃�0V6�5̄��n�{���D��`�|g���*���Vui��e]^��`����.v�.�� 8����~ma��u�gsxC�x�����?�[���D�0�q��K#m7���o��MU% ��%��c;� :�*�7㓹�!�M��S�KhB��r-��G���m�Q���Z(	|A���B�_�x�Ҟ=g�u=�w�~�q[p����e�A�I�d��(���]�f�3�#዗��y5b���|+6���	�`:��	����7�.ҎgD*� q�UZ�i���@6^��/y�Y#�Wrh���p
��.$�D�Yӽ�e����&����jʿ��>�@��T:]p�p_w-�k/��8�T ����7v��*op�ie���d#C�*j+J��\���̬qbg��{C��a�z��Y+ۆ�����W���_:����&I�.P��٠j�I#mi �5������u�W0(�즁������ S]F�u���aށ�P�7���M�2�fp��|v+i4T���_n7��,�%@1��4��~tRKe�U�8BX[��]�z�����`��W��:Tql�Yƽ�(vg4����/�=�,Z-��}�<�7?HDμ�ęn�]	{%����NT.�:>��n���
 �5W�Q�
X��1x��"m�tR�ޟNݗ^J��F��:%V�֬L���]d��Ɨph�-e�"�����BS�"�Є��e�ӌge9rd�R�ްY����c�@�񰥴@��(��x�/�9�S��uK�@� �V�����0����r�䨷�,��b��9��V�KGj�&M�; k��ޡ�܄5��4�L`y.�g������5�#�
��i�7���"���*M��̗�5�6g��UV����`��`��4���N:@�A��꥗
����H,��(�B�ep�.x��>����Q���< ���'�׊N��YM�B|. �k[*$-�^���!�ה_�T[w]���s	��J�ε�7�.lx� *`�	�o�͖y�2�r�(
n��߯�o���W fd�//���Z�>~ l�>���䡴o9#�{�JHƕK�b	`�b?=o�>����������ט�6�v�_�:$�.;��o<(�7�)�R[2GP�!�ve׮]��`v��Y��x:��?�fo�i��h�4�>;o�W����9�H� y�2)�ݣ�] ګ��]'qZ�A����g��7���nm�@��H{�.���ێ;]<$��
^��y
Ի���0=�ӧN�`w"6?����~���7a��Z�!�k��Am�knL`u6@��şf9�J�,�7S�P��L+3�N��  J��E��]�i�y��#����:�ېbd�eT�6�$L���W@�d~]���1�u�M$,փ���WL��R�>��� ��v
z3��ZT����� QkVT�6T$O���n��˂����N�(#"wVL�{S1(�y���P%�G�ȝz���=0m����rg&��_�TO�ih�ȟQ��@��:W�e �$O?l!��A�*��'��c��+&��n�=sb�.ŵ���:ŝ;�ԁ�
B/�M���-�͸���DV�\�>O�,s�Z��,,ۭ�.��V�������ǆ`5�~�^����?�
Em�w�}����Fl����V�twd00�#�-��	-o�2(��IfN=f���H���Wk���C��\U~æY� r�:�j2�Ж���QlBb�Í$����L�0��7��Of������f�����f]�%�z���Zɕ��F>z�����]��P�1ŬO�a�N^��S�4)��u���K#_Y4K�)u���8$�{�~	�Çm {�a�EDD�yx5/dc�j��V�1�?� �J�o���oM�;KD���2�t�? ��H��y��/`sh������b���U�c+hk��)t{&�NT��ei��5��%`�D�oq�Q>��	}b �L�%A�BEr+�s��sQ`B��oa��p/R���KirH!&�����CP���F�d}PC��,��[+�7��J����&���.AA���8�K,��]��,����A����cɂp���x�V�G��C�%��a���c3�-&�Q;�w|�<�s±�pl|�6�O��$b��>��d�U�����^�/�zN���������+��e��Xn�\�M��S񬷠�M���p/�h�]���|����Ӛ��91�?��ı��7��O&O����M��
�1��aU���y���s�c������nb��b�t��w��HUo�歼w;��I]���/;��eܾ]oZ���s�w�p�>�C���O�^�����o޴�CeO���n�d_�H�8�b�:?���V��-X��S�7@�%�>�M۞�ֱ�e.�m"�ᮈ/'3}F:M.�U`���R�gs�@�ۇV\�o}}�O��]-�4Oܳ;F��[�Ө�-Ļ7�iI�Z-!b�T�N���L��Ů����M5;Sz�t�C��e�">kF������?���P�����^0������s˳���1��ؽ��� A|��g���ބ�>(�z�d�V����t?�i�E0,�^�:��SQ�
�^A���Ù^���6��-=-�cm[�� �W=R��G.5QR%��ߛ <=2����k��s��m�j�M�}ὒشѿ¹vxx8�/���^ۺ�0xsySv9e1�5c�֓]���0oAb.S=<lH��ɢ�-��!������?@E���;/_�\{y�u�(��9��/Z&��T�t�=s�E�i3�q^�zzz���C �nO�.J0D~z;2��C�s4���[9�Gj�?�QV�k��"�Ж=jh�����w��WX��k�k�XBػ��6�K�XX�#��r鮲@Fҝ;w��lR?Dus�������NP���%w����VP@����JS���/D�ʱZM��I�#�t��8fM�%���j��0��1�+SQ�:�q麼���]����Ճm�ɔ�y�yU�"�L����'gm{}`=����:��< %!�s���2���9���51;�E�q�g�啾}��n�[���b���p�l�svt�6�J"��}*7���B�>D��Snl!��k�W����;�ֱ��7)��cK�G�����7�ƒ�H��*�!�~?@T7�ڦ\�򩄬��q��wY��6��yDj��M�{�tc؊���=$��� ����py�l�0>�%�ܜ�ajbR�Q�O��Du�������`���M*�"Xe-X�Ӽ���O}�����!��\m�xE��[�wL���gߒGFF�
̉G����$�J�MNN>�:[�Ј�߲^���c��?�-'d+���ӯV%7.���Lp_?y��R��q��Zi��g�
A��K�u��l>g��;���&�
!�\.oR/0Nj�1{��>	1����"!z8�&�.���mdT���D���L+�L�y.�;`P�]�m-荣�?~��v@*K�#L�v�)�w���I��7Щ���+B�g���Ͽ����YQ~�F��9�!��TW9��{����Ǉ���zk���\.�eO;�yYA��>#n�)3��v��V��{IO�5��JNuɱ��ȴ�e�+.+w�[�Vg������.f2��\���i����)�A������@�q|��u5������q��J�٥�	�s'tM��^��]�X#���7?���������I?Z�E��d���D�,��9[�O��A�%���F�Qä��ߩ���!��#��I��?ݹG~=`X��F�Q��4�����==�6!�k]��x7S`��u�VE+N^�VYuu��!��z�0-z�O��h�l��$�A���n�銻;�U�V���^��l0��u��]GZ��j�x��񔁡��C����'�7�o�8 @\ݓ> d�8��9ƉUF:��#�������7�5�A��U�&��[�Bg+�d��΃=�6$��@v7i{MQ�-8@�[G58b�_o��ؠu2vi��6�2W�X�Z�V���ӷg���L�!�˟n>N��j��O��>���h��J1G-��?u��ڮv�̔���q���;RK�d%�ٱ�x��lo����Z'5�F�`���w�h"�����^�¿�����3������mf}���3�q`�r1�����.('��D���FF!dϗ8��󙌜��u)V�B�~ġ�T�Z����q�1_pyjM#b���,���>D�9{��m]Y9�G��>fv����T��} s�i��{��AX-�hi-���������T0�%]�v���=�޵���&���WC���D8L���Ǐ���m!%�_se�����XTi��I��o���%EW�<�u�~�/�s�C���˿����U�X�����t�[� �nlkk��$*𤗖��â�;"K2u�m�s������V�� \�w0�&���������E�:Ւ�W�`
)jkL�ȣ��s�啊ʝ��?\����<DiUp�MÏ'j���]��'m�>}SM=���WR}�z~9}��ɍw+���i�E����c���W8s0�({�^� ��2M��A��
=z2�F�+�ܳo���Hɖ'���+y��XPD����@YY9��Nk��V�y]�@�1�+,�&ɔ/�N�?4I$4�5r��tχ���#C��d@�c��I�o�+��tA6�E�͇�� ֝* �v��z��w"�j��oj@�� �ͺ��Z 3�8�Z?*)������6���K��$��8Ć�>�����꟰����M�j�~>��9�<����Kpp���=w���a�N� �'����v?j7
W{<ٖ{�ں���q���Xn]ط�NI='�d�G��DqP��C��B2����!C!���2g,��%d��92��Z��y�������[���k�u��Z{�+A@�xR%��?�]�`u�ǘ
�7X$�d����
���O'�=�z��!����L:�؟�� gBJ'��qiw���h���q��0��}*ϐ�\�T��>�����P�ē�Z��Wl��w=�Y���G����������mov��D7:^k�p�>��&����۷������ g'r'w���eX��R����N��:	QS�l:g��W)C����bi�xV�;�E+��i�*�B���9�0�
�x׏���6��r<��A7
)�����d}���.��j0��������U2��z���7"��^pb2N�b[�����W��)3�p���V�W&�`�_@��	��S�����1�+���[��~�#��~��=,}���ӀN��4�Z�w��Bl������'�g�&���x��^�v6���#<ˊ�h����'��d��,TW�5�f�a�w�a���_ �5�lZ1}|����U��>`�Mr��)���! ����O�G�<�I�b����9F�%?^^�����67HE�����@��|V�f���M�z�� ��s�A�u�]?�gqq~]��`����}�n�$?������1��Q���[�n�h�+S\�Ad����f�hN�,|���	8��I�A���,9yd9$��">��/NVrF��9��,m��������M��"[~TLH���~b��k�#��J2�
(=.� �#k0���gr������f�<���H���F�ل0^��u�ͦ�j�,77W�d�/�$S�@:D�&��{EĆ�%��z�/���D������-!YVa�A���m`�Ǝ��n䔿��孉��ˀ{�U�KiԈſ�C�U�^�WX;���##�k��e�HfK�wm�/+�<9�'��I�&LD����֮g��c���Iɐ��ЀY��]���#i)�+�Y��,k�k{p![~Y�MI�"�-�0՟����O쑑)��kׇ1͕/V���%�L�x�p��8��o�."�z�࿻ �k�S��jp+��f�5��L�ԗ'�C�>�j���j����)h70<�[�Ա|ZQs��AR�{�to�WS)i���"E2&&&U�OL3��/�v~�3�"d�Q{%�՜��Z4GRu����ł�h�Jp*�3�#fN��m����
�	WI>T�ܝ����G��M^�65������Щ/ �a�k�s[����_�}3�Z,���b���˳
����5B����0A����}��C�i��]h�p�g�㲣]VD�vr��T�/9M�Y�'�J��zD��4�vPݿ�N���=��g��t�(���yyx ����/vPz����+����Ρ��l�,m�$�9w���?��*�Gs�Uh��HAof�U����?#;w��\[�r�ק���ι�M�"ۇ�&ơ�(����R�f����:m�r��־\Y���Z����&����MӦ��O�j�C�i)��z���f�A��}����4jPT�)��.0Okt �m���ѯ�|p/��!�|���
ܜ�WV-o�V%�j�YZckCC�=��I�_���|�m����&�r�=�C��p�Pb�"��vs�̝O,��~����S'a	?�A@X�죎E���/�=�?��T`�F���ԝH�3�#���y�?��1:�LW���}�	+��P@m�}�;9��=6��tkO����d�S�:�%A�ϫ��U����g)�pj���$�W�:��N����:D{!�q�P�=�i\T���3��������P�/�+VsA(W�څ��-<>�A���&������uB��o+G�7���z��=�G�9�0UHϱvEA1��zb�����N��^׽K"%`���>pްc@���٢�z�X�b�DD�\|���}(�C��D�/�m��`�ƪ"��W�����)Ym�F�>�A�r���Wp+����P{#�=��ǎ�kk�����}�/faz��5���v��!ٷĒ	ҕ�HZM/�/=6H)}c�Ƙ�B�$��_�`=�I�2x���e|��@R�y�_pu��ǖ�
UI�ohhK�z7�˅�1��JnZڠ=���E��n���ԕ{�/?9��#�*�	��N����<��2�T��&Ӏf ��x_�����h\����e���\ �q���N�5�b�q9��>1~�j��q�?�P��ZHW�<��o(�8z�Џ����Փx�B𢯯�,*�Ii�鑌�!$��k��W�\Gۀup�y���h\�X�/߾}��Y�JFk�~II�������R�VY=�Co���#�?O�f���Һ������:L^g!��H�%2G��?���ur5�RGW_3Ңq�"�k.Qg`|�x��umD����'/���f1z׾�U��]7���_3��H�p^;�,������\���NQ��m���d4UX����3 �"�lxx|��p����!��p||�K�˦'�4���
��)�R�T<���)��S�l*e`j,G{ڏ�'*�E����*ǯ� 'M�o��d�����ͽ�
�x:e[��X����{��b�~��$���f�{6�S��j�C���?v�B��,&Л������l����>�}q�S�D�\
P��,q×�#U��Hb0�/�!p�'I k#/�ՓA[\tֲ���Đ��D�~��������`);��2f���"�ի��J��{qe�R��Q���u`���lU�z��d�9�7�cY�(D���}��ڹZ4�pq�?�m�WJj�o��S+T|�u���vy�X�A����~���@�Q�|e***Y�����%�R��c�	o��T�~�z��C��,���"5A_�.!��Si����x�n�fi��X/��8+�����X���qn��R�Gaވ/zKhr�x�C5��q�uZ,��뙵lr���/;�܊�E
��,�߆q^mU.
YYUN�X&V(,��G)��n����+�J�e�r~�/�`�IQPbQ����~� Y�R�IF��	ׅ�Xb~�}�C�jw�n�6�.A��S�����Bʔ���@�_���ů�2z7Y���8�-sQz�A�a7��*������"u:�Id���O
�v��j��E�Y��^��� 9�?u����#�-��ªA1ovf��a�F�Vx�g�n��S�x⦖����Пl,���i>ߴB�MV'.�!)w�6�d+�����IX�����ԑzSJ# ���M�5�SX�||'�5l��NT+��db}�~�eF���˿���"�y��2�.��m��ͯ�ƀ�+�j�K��¦n�M=����b�f�����5Pߔ�
U���
���NcǾIi��Tj���Wǻ�3���ч���������W7B�� �R�%g E�Kv-��'y4CVc ٢/��r"=fi��:010�{�u��9j�oo.��cSʂ4�n\v_�6<<\�:掶�}�a bPhjj*�,4���R���ܛ=�<�1]��=z�g@���S��I�
��{�8�{q�5א�5-� ��}�S\��o�o�/	?--Ř�M�%%�Q���H�����0�B��"��ώ�������;����&WYBmw��P"��v��Wp@���8~	N��g:��D�ʗ�q�OW�Kv�.�7�%�l�x<�Zw�5��qU������v��n=F	
r�Վi���9I�'-���?��3JP��<�w���J��}e��gŨS̳��C�"���^'k3|L�M:�������h	[~��Ǧm�ݵ�F�%���� ݄`��������9���~�Z�oFne��<&&&�����zE+����r(M���i}��Z�g��CƓ�Ȉ`�����\��}`�M'?����j~��)&D�t��ӆ�_��D�q'�R������>؉���~��)���ȿ��~��R�O+Rw粣���=���?���B��9�<CZY��3f�� ��^����R2�[P"pj��ŒL$�}�A[��l#����b�����O�.�g�n����|�V�B�p��"��5R��r˔��&]ՠ"�N�/��}�'�"R��'�'�-����G��Y4�BD� Yw���)�'o�xE�]�O��v���]>��B�/V0�M\�'�2���������v4�v��:��mI�B$m9��R#�`�D���������Ќs+�#��?��
�W���R�ΐ�#��$�4�u�Lƣ�{���
x��/0��w�O�	{����-֣\,��>��˥��+�/yȼ>�i�����'k	�=�D8$�� �<��?2b
/� m5�jO<93���ۥ8�(U�/C"���C �%g�OC<�~�]�9��6��僫���mbA�|��l\\��ec9r��������d�1.C�ڪT?�G�#q����j����EX6�T���w�E�z�H��gj� )�|a�64�_�Ʊc�[����{^��O�I�e�Au3���9��eђ6���]���i��C"��	��ov���������ĉ����0@�/���9��X��*	"�P@��.���،��mJ>~�h@��V� S�~��-�]�#����+d»EП���F�ʛ�*�`r^u���2�췰8EۥZ3>�\� ȥ���p0ƿ�$���/^�5XBer �A��>,M{�V��]s(Y��`{/O��l����p���D�}����ܘ?�p�mP�٭T�� ��X
d��Z���P�2����P>�9Y{�!��y�M"W��Ī��n=�Erk����[3����}8�֨YW1hFqI%W��:zd	�O/'��}wV�Xl�D�	v�ky��Ƥ-�''�h��[T!���N>��8��T��@,�`-Ӈ�d����*!Z4��8q��vI�a���"�r��i������+�h v??�������'n���k�����W�g1B��U�D]�
���5_�}4
�&�(j�	.��oF�% ���7Q�D*�`��\s�N؁� 4�o�S:�y�?$ݬyn�T��Ȫrѯ��oԀ-Z�P�Cv��,�Q#�Շ��A2����ߓ��/;���`(��92�Ǔ���:����_2���r!M�W�ȟ�'�Jv������oEz�����<�ڸ�xb���---���:�A���O��K�Y�r7I�Ȅ
��η�9 ��Y��(D���$x� �u��^�C6��BpcS�(o�������i�ErN���j���/�}�ÎXˬ����NQ�%}�y�7i@��w_lC�!������m�ԝ��L�C�?7Q�$�M��w? �1��U���i�Z�O�flb�!	�����W��(,�\x���rk둶b�rϿ
�w._V���%�9�ޤ JMƳ ��)`<�#�����4"���M�Ż��?M�D�qƹ㦓oI>YĔ������6T�g�A��rL��0QG�1����@�~ʕ�@��t�d�`r�g.�&՚%Rճp�c⣷�w[��N�8P
�1#N�Kb43�dDD�qdR�N�J��o"T/�ju+|�G_�h�3K�	�Meo���̇�t����ӿ�M�����2%W\�W�%�l�o!{`
���Vm*��F�E��,��a{v�頵Dc�}����vL���x�OU��8	Nk
����W�ʝ�fiƓ�����2��E)�`L�X:^2|�lD*��a�v��w�~�B������L�&	��@���^�Uu��X�x�6�'�U�e�jPN-�cנѾHy�0��P�K�yNw�>�ڄw��꜁��nZ���PrX���4��	Ђ'j3�~������a��m� H�S���a3A%B
u�\]+������+�ݻ�S%���yZc�#�7͵�X����j&�����?u@Y[1|˧�<��jV7��d5����yŵ�:�p����VY=���Ո�wV����-�,�;B�|������ghu�I�kW���}� h��u�RGA�D0v���!))Wk�J��ܠ��U�A�i�k�ڋO>��?�K���kI'�=�-.���v�C���j���x��l�9�!����G=X%S��k���Q�����G�*�2�WT�D��>��n�U�����4�?���T��h��8I����Z/v
�Et��؞[�O�B]���/..އ-'���ߥN�E��[H����Vۏ\����t��> ���u$ٴs�h�Cd�y��'�`�T=�I4�Z��p-G�ip+A0�G�^�oZJ�I4H���%���X��,��;��K$p���Y�>0�̭]q��-oo�A`�Φ�x,�,��:y�ONS�Hlц/ҽu��������e��=�Ɋ�a�8���5�����c��:��79:	-�-��%���b[�|�]b���v7I�`��{�/�q�'�R)���������&�E�Y���:e�kk^0䛘a����	N��g�{j��1���[���~|����xx��뉈k�b���r������0~��_�_&��"�'7�;���-h�o������:��:�n9�S�[���_��C���}���:n�^ K�� ~�ۆB �C���VTD��O�TӮ"�X�\=R&��.6�:��&�i�+�
)�2~Ư*E/}Z����Z�&��u�Ux�5@yţ���o�_&pG�&�Pxx��@���@]��`k����sk	��|�j�Z
���ǇXɼfD����������]0/���$ԲӺ�3s����kؠn���Ǽ~�3�N�e{�����m��a;�t\�9_֚Yb-��hp.�S�X��4'V���y< ���;�y\��f�� z^��@����+�|�~� lF�������I��PXX�8I~ r�$%��,^�Yn�V�0Dsb�\\5�V���^�P��'s��Mh��-��W�!	l���^�,����-�۫������϶���g�4h����g	�`+��Z�@����D��;�v��yS�|xs���lњ�:�` ���6��SYYY����Q�-���.Q$�3.��x�g�b9���s`��F�oI���N�<���	�"��l�����t�����"�,�9�V*U�<��)�#^�'��2 eN��(�'O4�9���w?��]7�o�i���;E�G
���wp�2 ��g`�3�p�|8��R=f�1p9����2y���ר酸��0�<��B��|׆@�Ҁ�oI��O^?8��ԁ�6���_��2���Z�y�UJ��}׋���'6��ss�As��. )z�'�a7��l����r���DTl���x�!_J@k��c{�p�g+����x����
^<��h&���M�!/�>�`��������������ϊq��8����KG){?���0��� B�����L9l�6�����ː���s��ţ������f�F��}���t��Ej��Z�!��.�8�	�Yꚛ��FBq������B�Y�}>d������MB$�עiI$	�V&mݚS�t��N	��-�g��)���>�U�0�3�\�FS;��܈�����G��F1��ƊP�b����Z�ڍ�w,J�n�����V���d.Xf�Yy���䤧̀y��N|��'exI��6� ���g�>�w���P#�5#��0
g��d^;�n��G\��������
b�wq%/H�I���h�%�?�n��yL�L��_H�m��p ��m��!�as��N�p��|����y!�y���eMMMo�ƌ6X�i�D��
߼pߟ4XHkO�#`+w�3���`ӆ3����u�T�y�U75����m��;&��%[�J`���2��,5�-#�G��`�o�^Iޜ�����8�eJ�����R��D���������q�J�MUeew`2y66~D5膀�+Я�̃g^���v��>ò�J��!N�\�ܢĩ�̭��&���HQ���ލ������$�#:�\�U=c@��lւC�<��������'͡?w�ۣ�|w�QW����¦c��h����Z'�C�Q�O2On���0l��$�LS��5���/��թ�U~Z���C2%+� .�h}GXASb��n��H�K�&V�^>~�GGǬxO��$��c>;���� �czH5H޼�6ޛD�K��">
���%���Bo�H25��/+��^A^�>y�k�y��mvv��@k7�=d�
�&�r�ib~��R�F �O�D��]�ғ� ��e�@s�P&��Ģ���~iJ8^�������mƛv�W�^��w�2�D��UI�OL��Y퇻�o���ln2��0��������� !�$����+ �8���[U�nW�MR�Q�VV��w�
��"T���p��BZhH`Y{=���y�aGN:x3������&ĐΜ����*N^�%�(��rf(�3�(fIh��7YR�o!�0M��,�u,�i=�/��E�l�����?).�d��@;���'�i��%�������Z�k��1�w�h�B���mҞ��\%��l�?��M qȌ vpQoR���|de�^ԋ�9sbU�Γ(��E9OӺٙZF~�U��ׁ���߿�F���/h�����4���
�gX�W���$1�uݭW�澞��qxƼD*�ҥ��:��u�2��:��;��W��7���]�(�LD�}�c�����+�%������͜��Vŵ�1L_�=�J�h�ecFj�~,��~t�ݹ��ˎ�����ʃg�Z�k>|zy��q!��{x�\�Ĭ����Ȇ�j�@�y�������vhǽ�U�V��г�eG)����>魪�;���`�ׁ��R.��L�`�X��,�#�[�>.����B�QR��V]]M���b	��{ʪ��0����HPw���n�jx���@^O2�;x���{�k7?��#��g��%������Q�>x�h]l|�F�8Ԕ�^����N�k�qgf�VHp�]�'�<)�̬>Қ;�K�ACC�C�扩Gj=6#8	LO��v"~8{sx%�Q���{PU���;��)�Ma?��'��N��FX	H���.C�4�	Ss���;�4}����+(Y���Z7+�A�����/0������ZY��;�4o!��gw-�v�]
z����9�tH�;"Ov�,a�ٲ���������6�~�lo\���'���o��j$�����<����\��)�� ��f����.>�>v�M��)81Ծ��C[U��OW�C�Y#Ng7T�ՙ��F��3�l[���>����#^�T=��74T�����`p�����p[��oʡ���WGX88L�ad�
>jYV�l6jǎG(��w�u��F��>��  �xȑ�P�>Ԕ�d�ϗ����E�|��'��¾$S;/SF?㯡V����z�����ޘY������?v�&��'�^����{%�����W���]Ğ���#��V(�/�j,/��N�^�nY�\�u����b��^�nm+�k=^F�n[��|g����of������r��r�/+��E���FB�Z������MC���ƴ��*"�{ӆ�����[%m�5��sy�S=7e��+N��|;��H,�~�������xl2�lp�5.�sv5��M�O�z#L���59�&��(�<�~�ݑ������q�_�#{j�X��(�l�*����̮�e����-��ؕ7ݙ�pV�_����kXM�GݻwO1�B��m����%)�\�lV|8_�w���_䕏I���s��[����T ���o����e뺊���HN0��B�,Qw��_��a������1s���7]�z�񊲕#�.��?��C�>��D�M�R�-vN���a,Wsݦ8Fx���-�݆j.-�R�"C��U9������~�]2�E��ǈ�LL�H�ѧ��}���i��2�4�#���(��WQQq�.|`���Q���q�ĬW�2i:�Mg��j��l[K���b1��1�����ѼJ7�u]Mߕ��\�Tt��-|�C~�.�����gg��M)���������
��[%l�O�B���a�P֔�CN�L��c��.x֡V{e4��^���FMԚ�-�C��3�g`5�\��sqɂ!�n.���`@ۗ���K�/��N��l�x:�bƏ1=K�$9l��/ W�r���Tw�wH.e���ϡ�T�m֠������Ne�=�xt����:|��ޣ����ɳ,;�:ɪ���M�����EF}�1��Â��)�D��v;��$�X�������LVuZ\ͨA��2䨨i�C�/+�p/Ӑi����V�Ǎ�ljMsw��F|���+��-��s�%'bh�`@r�A��T˒�f1]����Nw͝���ˇQ��'�h�Vv�8�:r�o�!����H�6���.����>I�8�������*]��8���w94�*�.E]<FFb��( � gr�Hc�s��f:��"������w8�$TKC�?��,��f��1�i���܂p� !�;�X���;V�ׁ1���sn�b�:~���q��L�f	s�����62��_N�,�KV�?��֡��B��<i�/}WHTRI�hg�=�W���~�~�~_�@��S0R`YJQ��D�gyO{�E9����h��p�������"�rQ=�dG���_�0at�_�}z�����Mn�.��@uR)RF@����J®��S��db7�\kў[g%|"��ua~~��N���b7c�I�tU�G����&�E�����Z���I| @"�2���u0�S_Y�E�]���ٴ�����a���(���|A�r5�6���r���F}�b1��w����E{ى0e�>
���}I�O�v�vj�m����m�1h	�����Բ��?��fі���p�g�`�nff��/�����¢;�a�6�ք�V��7ׂ�}>i�?���ĝ�M�p�؞�A��;L�'�e�v�)#H�>Z���7�iu�veb 0� ElS)
'_�M�X8B��﵅jU�z\��3�&�� e�(��PN����
�+��Я�S�f^�Z���?��mdʺ
̒�b��������O�T:��"{��jj���#w�ү3{y���V9�5����Pϰ.�V�� ǇZ�~�j�G���5�، 0[��;���u�k�����j���M�X9�P�	 j��x=<'���o&�`�<�����R�4�M)��CGD�(�͆�*��
�:�4>��c�GǏ����>��|ט�˻��0�G������>�rգ��a����#N�z�~��mD�H��֣H��D�At��Y�X��V-��`���C�փW�U�� �������y��p�>�6l+���7$��{�&@J^���ħ)��9i�P++��k��BZ	>��j�O�= ^}�i㥈3U�A���e yA��q6o�r	�gN�
�S(����i�:���)�����*�ÊȘ�h�^&�1�s�zdC�"���(i����2�q�c�����q5� �؜I|�����e�����e�")�8��V�ЯN_q�2.�h=��^墍��g�G��)��c�eb�ూϦ�߀�<�kj�T��S�%?7�8<r�q5g���Ϧ_�W��5��hr�"�c���$��W�yt' L1�=�>�����ؠ\D��������o�6E\�K���[4�� [��Us�����b���c�D��i�A�	e�S>EX< &0˘�ĘyP8~mpE�����ٯۛ%r?A��>�u����m��w큔ѻ�Ad�5A�F_0/��x�Ӿ6�
�L)�@����v��
"ux9�vƞ������K.�����.]_���jY���JLvJ��*��|c*-�D?�/&�n��q�E	�8|�:�u���4�pK7�.U�"sQ�PZ�P�7�"�Y��?�oW���]Yb8��+O�rl[+`B}Ssq*E|ضH��ӝ&q;;0�P���'Z�2$�'!aB>��2T�5��&�����U%�;M���߭W6~,��{�v��|�+[�\�Ӭ�,ZQ�r��d��˷�(4�[����~���@͆���Y�~��x�/0�����ö���B �q���JH�A(��3�X�G��[?�|��,e���CO���t��a�`U��o��D/�����
X:�ġuBZ���gr���ޅVK��É�]�!8� v����죪!������.j'�a��6�J�4���!���늚h�F�����V������|�k*)9����i�~d*��z\��tV���&
�gi/M�׋m%��u&�ieW�� 	�k\�M�}X��*+G�CC��fE��\J���i�tqll��>��l��X&��#�M����N����n�]`��&.�i��:�F6��=�aq�`(� ����<n�`�RB���Ԝ�#�M7ɷ���s�|ku�o��_��� * v��ady��ի�K�奁���P\o,C$��8w���M7�	�e4��h���T�,��{/?�x=De���x��={'��
���*_/�_D�������^�$;�5᚛�U?���q�k���|� �7S0_i�M��r|m�'��n��ی8|��v!�lv�6�'��+%(iu&&2����;����+��#|���:�72�1�惼��!��6~��C��-[bˏ+��_U�	 ��� �餴N�49�pLr)�U���G������>j�/����ߨ�`������~�q|���#G�(^�?
~t�� ���ھM`p��0a�L�_:��U�i��i���7�F�L���#���!����և�ԨMa'�݂5Ƹ+�r�U�/�ؘ<�� �f5�,Z{Yp��P�P�|��&�
�9�ǩ^<Ŕp����G�JSJ�&��9�2Lp�p�M��Ʃʪ*C�R/�+���h�H�6nʰ^��Ǯ9�W���{I�(��i���t�Ѷ�hz0���P��W�[���<;`�𙷂|]�,	�~����.�5g�2�5��P���h_���n1>�|��� `�W�����J�qW�	�#�3??�n6�)��
�Crc�b<l�CvK}�~��Q;�0�H�t,xʏ���ه�.�M)�(��g����n���$�֘��/S���X@(577��HU3�#����	��l߄�5 �9�O�[��|�R���' ��������f�ܺ7a�� �
 ���Sǔ������+�n���FpƏ�V}��KA��荫r�1u�y���m�*ii�	�R�����a!�3l��2	D0>n|R`������Ν��W�:�ດV�������&�Y~���2<�\ĳ�4�3���� �as����p����9��f<�0q�����VxI��v�Q���?A($�x�'��94M5E���S��Ņ��^r*���ы�:*����Egps����u�@���!Q�ᆻ���eg)P�,uC,��"J���)�w/�߾um�O���G���jcZݟ�^&l�����1Q���*J>�F��T(�r�ۯ���m������=t�	x	S��W�o�`�8_��Eķ��;[Y߂��^�MEӦ��� ʘ���O�1k+�X���=>�hB{Z^t7�����gWs����Ǌ/��#��3C��CY�I�#���Sy�V�M�6�_K%����'y��5�f��۰�)�a!2�2	'ky����[��t���8�]���X���H�n�M�+yY���R����>\QQ���L�+{A/���<A7��/�*��/�^�;qiiqa�hl�.�w|$�2�d�ˣq��p)�JD�!�<����L���5�����/,@>�n��*ڳ���qż���_B�[3>�ؐ�K�˴����tt�����u�#�o�b;�a�`q���M���O�-X6l�i�r�3�~n(#+UWUҊ#��u������X
8�""�Nоb^5Q|:���V�eZ]��M#G�y>�9 ���GE�o��a)m'�c��cX5����-�c!��Nq���Dy�I��t�ޅÃ\	�� 	�}G�g��dAn �s �8�ƺ���L+`L��]�j��PjM%��ĥn.�_I<��Ue�NZ�&&��IX��3�Y:2k�+���Ha��S�'X�h�� 8F]�gS\�p��q���P[h[P�����Y��[��,�8�O�.��]�Q	P�Е: B?�a�-�N)����5
FO���t1����ծ�4 l��? ��)(>�)�"/ʷ�"�m�~�=<*jɏ��/9uV� ����n�*�6?�-�oct��݋mv9��U0���2e�<Ho�X.������!Al���q�F׻D�+D�Z$zp�$�	`�U x�qc
�]��� �mA,(��aGj-���NFԏ]�kY���v�Z<ʬ�/�!L������I���X\y%vL.&ڟ���wnr�͈&���?<`8ܚ;W�Zp�)˾�3��4Fٱ���	��]�b �������w����[���H�<&�3�Vg��Q�oBM�����	�r�����Q=7��<熰#j�1�l.VA�+:��XC��.���,����㊡s해�ʺ��^{ѯ�����j�f�¸cd��s�!�p�����S;v��y>�*��<�������Ç�<_����绐});_�T�B�ی�W�3��ʞ{Z�*<��u?��W������ RC��+je��j�I4��U�|sd�}G-���{�yx�џ���m
2X�M�I��*|\��p�}�">�mJA_EN�%°��zsG����X�(|���	8��ESim�z6�5X�?~ �x��H�	�h��`�Ƣ��F*�~{�='�8+&��׻�I���L��Wӗ�	�Z��8����;�n���D�0����(�$F�m>��ӄT��V�����+�l�.c=�\W���݋*�g`j>�w(�װ���hϚ#�����cT��Df�S�/,D��
�X`�"�*x���tDR��� �V���=:�梇]�F�>���aw�v�2�#b0�-�5mޞt��D�vt���6�ߔG���* G�j̰nӭ���oZ�w�����q�M�����L�q�6 �K2�]����XW��\�A�V��hʕƽ�t_ y�uoc�ꝇK,�09<�*P�d�S�&U`z����i�LH������lp�8�������#I��Ċu�/��
a�BT��O;���8�¹�*{���|���rd ,���	9l�EH�|֞����-�9_��T�<s�XMMĆl8\��l�SoI�6rdP�n��*hᡀ ��v�Lh[K��\��	��1�0�|G���2�]埜 ����\Βd��L%k.:��߀�h��MBB{���C������v��6���Td��$��z�]6��9)�� R�-�J�~\auU.�b[�ǚ�i�Z�rL�g�P$�\��`�awk�qv�o�;���<�_�v��=����D�W}7O��l/�:w�[���y�e0s0�(�Ѥy���H�,�S�N���U�f�Ȯ0+�_�8qcچD	��=�i�A���hχs8��{wI�an����("X��qs;�pO2����4�h
��bBڣ��a?8]�)!�w����NV���R���6R ~�)�P�����L{-�����Dw`����@�d�fn��#+}=��¯����װ���涚��������[��o��4`��:l�E{�)�2u�L��\�@XF����ͨ����v���L%c�
������4�ه���3|��&y%?WU%׹I�L��òC?(�m`��Z�������*El �
4i�}k�u�oba�[�b�8R=O��`��U�!#�[/;�1�-!�Wq�K��!���a&��d:���g�@�R��<�j�i����b���Ķ8�a>�=OeG��]��\�������	�Fhh��f96�٧�P�ſ)��_3Y�r��4�WLU$$$�`VK奫RT�3��(���}�n�%'	9p�]��9�H��7
"+�����إ�ļ�f#ѻ�`��iE�R�G9yAEQ��񌦅�� ���-�)�� ������'�tu�:���YGi���a�ػKLl���4���[X����-���c�G����v�%�!�<;\�rj�
"�3�E{(�b͹Z�]��a2�%>Tb��w��	���7F�-ڹ��v���#�`��lmG��ȡ����^��u��?�9�]��XڇϺ��3Q.*ĵ&�,ż���:~�1]i�AM4@����H������v����2��;$Ꚋ��촷ogo0x �m����a�@��0c46ُ�_�C������B׍d�nC��M�wsIt��ٺj3}�M�a���Y�����{�6�,�Ȋ�gOL�!��1'�a�l-�9W5t�=����5���P�f�O���u˄߫������k�ҳP'��9+X�y�M��)��@��*���l}��{2�� �!𚚄;%��"�"�I�аx�K\k�`�����9]��Y`��xl'�p����>y���(���ጝ����Sڢ@vgMw��S;��{ݾ-.�	�� �\�����D�b�����6�����~�mZ[f{����#�%D�Qi֭���?}�?�Y��P�	G�<m�7K��Ad�ǆx�PW��T0A���h��P^
���/�b����_.}V�C�j�����-�*t�F_�G5���B�<�p�R��zN`�Ġ��ϼ��Q(�G������X�]���{�6䈝^a>��Aw�)�j��SL�;����U?��d3���z� >�.)�
�8��gp-��g0N�:����)u�Y��yFN�|/��9l�dC;���t����=pb��2�D��"`F@%df�����uhi=ў�Ϧ���@2O�=�q�6�K�(���{�������|ɽ��<�Y��j�-ķ+iu����@��i,b�J��#ys�X��gw���H�rɧb������
��v.�k>���Ν9r���e�U�D;��k���g\�/�2Y@֦@�E̤���t��BCV�/7sX����Ut6$����yG���5Ӆ;��Q������qH�v8f+�S�����)N��K��c>���l"?~�o�?���{/Ab�ݬ��bO\+�T��f�b�h���d-N�����}�.������������__�����k�&RF�	�L2`�w�f��}VN����W�~�i�L�q�C�tut<%���@.�L�����m/g���m#Q
�^S+���a��즡E+�i��������OϪ�=)��p�&�#L��W,�<YKJ�=���_��V���'��ژ�Q�~ɇ�������Ϸ2��$�H��8������ `a�V�,�M�r�J�k}�H�W�1�El���+�1K�5V�pa�����Ao��R����p;'�,ړ���g��@�:�{8��9�n�2��z|0�����(��d�DEY�C�-�.¼K������.�a�i�f����3�W[���N�����ܔ�`ç'.c=w����)|E>I��-r�6C�@Jʡ0~�a�6��-�����Q)�Iɽk.ߜ��E�3ρ��a�}�j/(��CF�K��o��r�
��*4��\F��q!cG �q\|���O�p��]��?Ɔ,5L��d'�,�rn�����|k� �fk�� ik�O��b<M��oS|��>�رwS���i
.��u\|�u�mV��(�+pd3�������6��K�j�_�d{&�Yp�&����΃[�olNw�a�<���f?�v{ج�ɔi6���qў�5���U�~/�����f�.v:=g:�'J�;���tԑ ���g,-��f��i4Z\�l���L��]�����Z���oy�K��
L�i9&�Ŗ�Rډi���.�!x��^>Zt{������\FeU��y翌��ۿ���oS�}��� ���V)Z�X�]���ܔ�m:M����fD����r�iΒ,�Gt�4��ǐK����r�s.Rt�m�X�N���;��CQ��zB�1����P������ND{&^t�D]��9�oX��>PgAǰV�1aB�v����������3����x�f���J�DJ�g��9���1]266f��.%�m$�7�E�Q�MåP�� ��ӿ`������	I�%\�6f�h��x)�ZK��H���W�#4yr������Ct�b�C�%��10����$w� Y�%(��ə��9����/d�4���NYW�����Ju�u��1���\?
v��4 cI���Q����{l��3�Y�,J4ў~�x,E)E�hU�x�#���"�[�9f0֠��"�R]��`�[�Uc�fl;Qf�8�qQ�-��I���h2g�_�ԯ�
(�O�����!s�#��0!9@��,�ȜRJ����+o3"`��/C���?B��x��>/�o�O��$�)i����/#Sge8�uW������t�=́�Id��[�&��\w�4\KY
kYVm�a�wa(�4�J$�7��Ƥ�ٷiii#�����.��F��$��2�g�GL� |i��j�d�S ���[�s��S�B�J)��$y�7��ucfU�g~�%�^�̂���
����^;��!�7��,�%i�}X���.ů�����-Xt1[RFG����4�����C���KZ1�F��VH��gff�۰�l��5D�# �+�ITl&��ؑ���^��m�/�CƦa�eo���"�Θ�`�);k�ӧݰJ��ڲHe�}�,�)Q ��ֺ��@��"�Z@D�@4k�����q��c[U��a��#��pw(�����4�|���+]E�(���q<�������	�\/�Xw����ᇶI�Rp��@
��>t��EZ��Hk�o�懐\6:4Yf,�0�O9r(��Nݑ��|�wh�C�j{Fr��6����/u�>��"ND��&#�ã	�C9�f�E;�f�jS��:��� }�������C�Q}H�k?�]���ѓ��B(هh�g�ډى����W0 ��bu��_M����-�nK�D�v�^X�VwB]l2D��YVp2d���	�S�	i��Y>�s9E�4�>,�M� �s@��k�z�&�3�&�%�	����&jsZݗ�+�aX[KH����T����EMb�Ђ�k���BQd�Ï�U)�MEv��Ԕ[�i�eO��J��+�-"�µ�I�e���s{������}=_��y��8��y.��RC��K�ݯ��ܹ~�_d�;m��9�'xg)������Sw�����i3O��>Ӏ��dX<c?�� ���,n}�����F_�1ڱ������1�,j����O������ĭ����Zȟ�� `�Wb��7 @L*�+Zb���4����Ԃ��q]7� <�?~Ïk�{s�MEI�/��1eOB�ƫ���c�\�[w�
񚰮YINM�uq����ڱ��$�ؼp��Ɨ���}��T�SǟN��iM��m���'D�������~�4_\>��USU�4���H�U��(8���%\�X	̚Y�X9��,� F��,5A/��on�l~%�z;�2�j����p����y��\�<)�w����|p��X�g�c����{� Uڸ����/=��M<�"D2���7��Ԁ��H ����: �;�]L��:�g)"�]�U7��B6!�c2LU㪳!�t�8Bw���%A;w�� W�3��O�`�+S�p� �����7	�	m_��.n�$��kݥ�6l���t]H*���L�a��
�x���"��XS�;|E��}���8%l�9[��hFaz��9F1.�Yyq���\UX���a*y�K���IcR펍���|��a�2����cC�ƶKr�f�!��1;�=�TE�b��N�B��yY\�o�j;(4Cq���ٲ
%I��&�����u ^�G�(�:�ښ!��1n
T�$�a�#.�a�SBB�p7n��%��{�j�K����?�6W�����ڲ��!���&J����I��tQ��'S��B�X#?w@�+k�z���BF��e[�M���M�E۞V�ꕵ�苩7��4�����Ma��q�`�����h�M�5"��9*��Fǯ�eeM��i#��
�^�80�0��`��N�����YQ�T����wBǊ��57"`��+*|}�S�(n ��t��Ь���5g2������&\�h�S�ri�"�\<��8��3�ρ��*4K��N���ySq�,��Ω������jV��>�р�
�A�9T�sϘ����� rp�+��0S�Ԗ�66F��E���=@�j1�e����	9��3��;   z�/wi��Ϳ���˃���0䝳���A���n���It ���5����Q4���Xu��E,�5��'�' �ZƏ�����}M�{�B�dP;�+r��w��Į�Z�a����f ���Zդ^��!����ᩓ5�����~�_�CKr��f;u6-~�����Rx�)<6��eq�:��ؽZ���#�]�L�М~�B�o9\K7�cՄ���;�����{���#_��q�O]�X�����-8�IղKLJe2�tara�"i�ם�f$��88�\h2�*�3��l�D�����m�[�\�I��7a_��y��9~=`�x�}�4:UZ@y	�
�\�q���V��KgXS����N�H����+�̨`�з��;0�~�755��wǽ����D�'�5���?�%s��O:G�AΊ}e��y���K~sA���1�Jw�Ahf*N�d3"-g?�r�?#��@p|=���4��(�c��B������,���Z~:s���&��ZgS���ťծ�p��߼ySa�
hH�ѐ&I�׫m�O� |�.�7���
cȯ.��p��[�]���
9@�[:#+��O�m�Cx��M�,��:
(J3h}�@��G�'������"�������)o0��m��� �Ơ"�iގ8��QD�$�C�l"��}h��dxj+c,�Z��&@\�|���1[f���d�y_�����P�K�u���6o��WT�v�{�]�������'�(��:�(2���E�� a��߷b=z��c��B��r�&QZ��름k�~hRrt��Zl/\D[�}�ɶ?Ο�[E+ڿ���I�5�g,U/���V��+R.p������K��|=�|(���%P撟�k!٤�yc���������������O\�Ӻ���b)�2N��t�H��pw+�Z�y��;GW�qp�*qa�W�z'�SrGvC��V[h�� �K�'��tuu��K_A"g�+&��?D~���3���טli3d����b6"zO�t)I��j�?4��6qJ�a��h��}k��V�u�������`P��黬!os��mO�#B\QzzG�"~�F����󙌫��<����C�Z�������H�">
�
^�lw.r/n���� �=��$ڟ�^�_
(,!����Ƽv`'WXF�9�����W��Ĝ��6(���_��u�$_ݵ�4\ס~�-�/1Ʊ�A�{ᑋY��Հ1��S�O��QS�A*��*�_ &8����n�
z	��B�hDhv�Yy�=}��rh�a�O�R��ttå�B��~$3��1qq�u�E8my?⸨���Im^���`�n'�@�촁�+�-6FQ��H}wO�3���t��b=�;t��ߝ ����:�v�v���Ut!v!���&�;cB�b�����5����������W^
�| FQ#A�YF+L�"�_@�h��$��j �<�W�{zyO��}}�7����JqW��8@�+�/�.��a��c���w;*2T[ʹ���u�=e��s���G����$v�`���s���A�ޮ
�sF��r"�*\TlR�<FY��|%�D`�����z�	xЛ0��d��X� �G�C�>e��}�� ��_��[xT�j�h)S� � 
Yl�/��rJSS����]�6]{Hdֲ=�5 *Q�!�p�q�6�m��o'2y���q���|Uە��꾝�ksN�0��n����صGNn��k�+�9�P˟`��3�V�i.؅�l��m�+g2p�k�O�BD�)��xp�8j]bNYO�������khh؝!�R,�BVQU5w;i����G�4�`�W�]�[�\��vyD�P�.�ͽ1�8֥��j��_&����|Ԁ�M�%p���{����Ԓٌ�l��`��/�)EҷM?g/������L~8�)I�Pm0)����b�3�ϧ�=��K��2CCh�)f�a��')2�MARQB.��w�ͬ��`]g���6��-3�Op�y�U9���Ou�}��L�5�[j�-���!E����"%��p�#�����Xvj"�;?��[�ȼ�+GpA����}��>+��5F�r�r����Td��e�;�ՠ�
��F��e{~�6һ�DPRw�jɄ���ԅ,�O�!h��(�5�n�C*.I8yg*8w��m��=0���T� �!j�@G��*��	V�C��ܪ���t���۔�N��H�
nܸ#�SFz�Y\�z��	ͤ�곴�%r�! �[╕�j׷����.*�z޾ p�9��ggM���<��n��ҢX�	j��.?����}�1��=���HNN��.�C[�x{�%[,�E�BW�N��:<��4�z��`aI��b�%�dP����:nf2{�Z�a婿[h��H[�� Z?�C��{��m
��Ox&��p��&�`�Bʅ �[vY�����Y��Z������=�\�&DL�E�t��.�q5�7��/���A~�ߡ;U@��(o�"@�,�ﴛ3(7��b$^��Xv��0z��|9H�˞�����aa���_�m>���&�0������]z��WɌ0��J�k g5I�M��Hm��[�鍐.�s* �ˈ�_%4�.H�,�K�C��H&��@M��;�	y�=[oҩ���'_�.K5��ג*d2���>��ٱ����L��#͑��D�丠�v�^"m\$H����ԉM�	�-:�@��|I�Kl�=�sir��0|�C��/j��AW�R��΅Ƞ;����8�=��t�D���g���l�Tܿđ\p"S�{�,.?�C����[�E��]M��NstL���o �VS�]R����1W�V��f��7���(�a��ꒋx���}��m�Uo� ?У��ǜ�1:>~��y�l:���<����:B�6VVVr
�a��S,da��e�Ux2���`�B@Ξ�g�?�	u�rh|���:o�vl��@��W�9�6�j(��BW�t���<xo%Ze��@v|Ι)���m�������rkH�Wy]~{���K��Wқ�}k�Z��S�T��t\Ѡ��p#i�J�_��ȹݽ��w��b\)"��M�g�P�^8��S�hK
(\��cɁ{GRw��\z��=���!�c��������n��b��2��8��6%��H�,:5���H[��-��1��U+����@-�8�;�ї��wR�������X�X�~�4
�<��\w��Ţ�`����zcV[i{���*\oӳg�.k/&��0��Z���q�]��=��g��yά�灓zc�o�\'+O<�l�J\��%�ң��<J?�Kd\��n|
�Ӫk� ��</�_�����!B�����wkD�+w��ʑ��Ǉ�X��S�g���}3L�D�ThJ��S�#��,�d���a��+�H��M
U1�:5��+7 ܙ����g����y :���X�p@U�R�L�_�]ۮ�3���6+� :�0+�Ӱ�]�;�3��&a��5Y�9�i��ͭ��������1|�7o޼�+y�E�ݨ\m����wa���;�����~�xZ����G[ɢwi�Ϥr�K�̮#��6*s9�!E���`��9�ӽ�j�T��M���H�"���Աy	�BD�p�e�;̶CD��q� j�z�XZ��>��G��q���}x:.�����Z�e�_�$.��o�Iu��ڝC�:��8����´w� a3�)W�o p[k3�l��]�&p:�2�i"�`�#���._ %��$�}G��$9�q�wAy���u��T�2���>|�DKCp�U�{��5�f��KO�ڈ�
����Hc�`}�;�ru<ޣ�g��v�;$$�7{ y$��A*�ޥcq|��uPR�l��=q�С%��,��pz'F�f6oI7l���G���*M^y#	����ŏN����/�9$�8�-���Z����5��G}�4=Ԭ�[�o�qo���f �-C�?/tI������q�����|<2�ǔ«!N,L/��x������cƖ��������,hb�d�?rUk@���^ rW�C��(c%1��V�*O���zx`��U�.��34o���M ��9` ���[t�vA��X�uy�"#��&��0z~� �&&&�1�=�� km�8�#`Dox���u�{C0U�Jð�Icu���Z�����v��[��92�~֔�x�F�[r�*q�,<��-��	Zz�r\;c��?|)A���-���t%F���r��W6~��W��D7���t�,�'�qǜM)}�u��)Y �z/P��v����\�.�@�u�MZ���9橞�d�r�~�ܤc+uϦU��	�������[IrC�������=����hw�\��_entj"J,!����U�Z�	��*�"K��4Q�4S����
�c�W�
���A	�/-"�!��"1�i]��5�\��h�ϻ�mC�뚥�e�q�mlZ�QZ�5U����Ss¶�����O_ ��]Z���ݩy�5�(�x+DN�#!X�ƪ��7]�^�����W/�J��+2��-6���˷whh����*�#���z��+�B$���;`̱�%R� ӑ'B�bmN㼞�����ih�˺��<�fP4�����M�;��
���A�?���f�%�D��#�"�����	�3 Lԙk��K������Ca��a��;i?�Z�$[�EdT�w�{���C���Sj?�.�j ��fB�����	���Q]mM��k���eaM���]@?�9;��q,�����R�= �u�#\eIO��7fgu �+��FЎ�?>�ϲ���NOK-�ҵg:t�o#�a���d�f�};�<^)��'i��Zn�!cma7��n&���KC������U�{փ�oxΠ��H�|�U�]zwO6��]�����%��s\��z�J���۳��0xď���	�����ަ=�RC��@.�Y�ibb2�=Dg�;� |����Z�5Li*��ڔ��I��֯&�Sn�8cC�eh����c���Kᙤ�f�ɒ���?�����&���K���C���`@^��*<�4d5�!��L��ܢ[�Kj�s:w��W�ܝɇ56����������ռ��"9�r�$s^��s����f�~j�q����
	��4���0+���b�-4]�����/��$v�J>oY�!��@��e{�C�q�p�������g���)���Zڒ[n�E6���L��_�5M�u<6xc*Ʒ6�g����:�58--0-�Ub��^š�R7��"�㌗��G����Ɩ��i����K��.͹�x
SM��C�I4X�g�)��ɬ��7nv宒w)���L�6X-믎��IvD�,/�5Dw���TR�k�yD�ʘ�O5��픷k����Z�0dw�4��8*wFe��.#��o���Bu�L������RI�2y����{��Vk�P�6�����0~���_^v�IT�v�3���Ů�7��<ؼv:r�#�g��b���q�N0�3����#��f�z�syv�y'�h+<�,�SG,����/�tq�����˵�fU�<ciU����0�+ �|������,#-��;���9r�t��#��*@Шn*q���
���zĈ�=rK�(��V�+�(/�����v%g �����7y/Z�����M���r�.�G~Nڱxx�����E?&s��_��z9w�r��@�Kh#>>&�D���M"1�X�n�^���h�A"���pQapo# ��} �vu(V�k���wv
����O*5CXgX�����w�I�j^�5(�"6\tq�`2��o�/]駌��rj���$��w�ET�Q��u����ٱ^Uٞ h��&��7]N
���x�����0�-�+9��,շ��f���`��Ku�b��"_`v������1�
3�? �e��@���8B��P8��(EB^�-+��#:x�:ٞ0�}`��oU�ǉsVC���۪++����>L.,Ց������f|h��;���Ju��LJ�p;طN1��d��Ln��Ƶ_�v�c��@<���11�p�7Xݑ���_�Å��׉6���$o�mK����o0��XR�Wq�;��umY�x�%���L�9�����X��r�A-��|}i&
{�P~Jh%�z8�!�q���!����D׶�c�^k�mi� v6TV�B�����cX�'</�t�y��\w�mu�"2��2~I�r����� ���C8�J^��1�p�2t�Q;qMS �|��u�:$:�3���pSY,u�܋�>��L�i֣ȝ	jj���9�C,��_BBB��v���K��'��{�v������J4t7�ӟ��{��)b��)��#�� E��[�t�`�ՋՄ�.[VJTн��"D������S��?�n��ƣw�C���/��X��J�T�t�[�d���l�� і��^+ypƋ����s�AC����=l^|*��P؝�l����F�LF  �Z�)n�"<y�3�ۂx޺��zB�ڣgjb��sF��I��~��徱f���-����m��I�f�KS���Q�yt����:�Y��Đ����_�S�J/�������жO~�m�D���,�;�L��U��9�D���8�Gi���G�$b�w��#[��65��4�Yex�"������lI����
3��(������+9%�v��
��Uon�1{a�M�'3z�쒷u��'Ak�i<��c��Ќ���>(�!����:��ǟ���(z�*xa||���4�g���\�����:D<v�$��:����PF�(d�
�����&�u��U���ӵ�5{����[l�o�ĵ�le�i������9�M��y����g�ɟܓ��sIwQ�t��4� H��Xj^/a��f�A>��z��V{qhyia����{�Ɋ��P�栰���ٮ�U\®����a	��~��d����'��R�υG�m۶@�� o[��	<�)�6p^)&�/�8i��Ka�!�Z3��$�O2�Ļ`O0*

�p��:�����\��,m�G�yn��y6�3����Ej����-Iy�%��#�pFϥ��03�b˚څȢR.�b�=C���^����
2��D�.�m+������
�n*R�����
�b.�uu�����%�p�X���3�������`CS{ǋ{�6���~1��ӱ�b�r�Z��$���^�1�����b�J4�S�&� �h�*����SI�'�מI-��U5�,c�߹�mר �����P'�8�Gq<A����m0��1ƭ!&c&4r���(�ͧ�C�qX���(������!�����ab�h
����xd�*�3����d�`q��}���b38�$}�&�L[w䅩*�}�0�.�3�'�*�_�b�b���c��7b��9��H��}���^h�@�a�2Ĥռ�Q��I'!�d�N�{�K�/��2�"}�U�D-W�N<�{J��O�=Eyܡ���<eB�uhI�mA�0y�:����ߛ[�V��|�@+s��z��[��"j�"rD�p��e�/����ix��+�-����	����)}{q�?� OSST�1���0�4�'����\l��R��Jg�z��j"�0��˵��B�c���f:�Z�8]Q��\M�왝]ߪU@�6��(.�OVWS%��S��Qg��J��?�m�ݚ�f�/ҟW�=�罌��=l����:X�����ve���j�!2���|�&n��C�i��3 �#�w�:p�?����(.�p9&r���=J��	���2�������m	�0!��˱���{�2!��C���+G��(�e��M��N����N	�7?�h�s<gY[���F�80�&�B�;��~Z=$=GAY#�î_��/#J�R��o��[�,��+�u�]m/q�c
���%ݶ{��s"���ډ�Վ����]<Vi�SU�o/ �U����q�ni"��*��ǌ�j�Ζ�o>�Ù�E-�����v�����/_���8�s���+��? (AۮG��&|d�$�H&'KP�L�G�1ׅS�Ґ@%���b���P���:3Y:Q���`jf��>(��Y�Ϛ:�%)��

��B?!�)��[ �)��k�!T�^{���i,z��7�1�����*�X��v��.�a�:��==�:��튣�3CM�K�6ѭ7��ѕ���c���[:=6t^ii,�V �\F/`P����]�q�v�A�8�Omy�ޟ*���g�n�r{{{��2D��;wdR�-��G3M~�[��I��ן0R�xH��^����,z�}Wo�Y�X4�h�o�4]�W�x�3��d�xP-����z�c������*~�X���0L\9���d���q�Մ�K��`U�̍!୭����Hc/q��B�(��8�Wr�������������D�1����hǃo����H�L�t�l�a��G`5��ngˬ���-@a벦�R����������j��$�k���w߾�Cd��x�Ӻ�C�����h��G(}��ޝ��R����:� P��v�B���v��)}�q����ݾ��zy�����%��j�u���9>c/��J}vS���G���{�dr�Ԁ���x��M�BZ-���V�J�/���jB^��ʁd�ŴD�^�b^�I�����j��g�RB3�s=�5�#�fya%����aR��M���\�&-��������?�<r�R?!(t�Bw�#uO�Y���K� M���&�Ů1�fVS޳,�J����ޖ� ����8`fN�=�� : -׆n�/ �y���?��(�(���_���{t� ��;�^�b�<	�x��!�$��,��TF�튧��������B� �^��Ԝ�;3����� �!�d��2ģ��㪼�"�?�H��}x}]d�Gy��Y�I��\m�H�@a�u娈�u6�|bf����M�n[�x�#�҂�!�I�6נ�9 �0�n�,!�yJ�\5�N��`E�0��WL��ů�G@4��F���k��E��̿j�VaGH6�7�b_.^P���k�w�<�n���{h��o4�%%�r��ʑ��%D�sV��2�8�X�!Z���IP'�n�+C�Hs�e���"X+=��S�� d0�M%����7����[H�����H�;Q��3V��������]���~az�,�0y^.;���F+?�r�i���i�|��\��Y;�P�H���-/�R��@�z0&zsZx������|�n5�20|.�����ʗ����TM�����_Z��z�A7iK���{�6���ߴ�#B�ȼ��m�_�rō$��U&?�M��	��֖t�|��R>D�=��u8��4��>Ы��6��I�Wӂ:��/���o��qx�_�Vh�\�V!�L�yU��K�$9��
�5��_��q���B_�Z������[3$�?~��$/_���Ro��Й��I���.���������)��Fȯu�+�=Z�7�C��*s�~wh�ވc�,rcFF��-:V��ϰ���>O�~ᩔ��a:��5zz� ��/�]OY��z3�h˒���㏑��_Ss��	!B�S�s�-ܩOU���o������5�=���{������N��|�O-�������
l E����
(Nj��~���6cc��=L����43=ʱu�֍B(�?�π�'�Lz@V8c�^8�/_m�������5A> ��g}�Ȳ�
�j��eE85��aM��=�Q��݀���� ����-�4�H׻��|,B����m$�o�H��)�s%��G��U�� �+�kJ���:褷3�矿��Q�Ǒ?~x��:����)}.�c牋nxp���N�@�ͨh�a�o�Tÿx,�7�>���7��� ěo˵��E�/���Evvv���=�^�JއE��!`��|k'�X� v�%jA���S���P�AC��3�e��x�Y���d�Bj�o�N����;e����T���r�������V�Ic�`/�d����ݖ��P�.���)~�]W\^��ۆWq�a����ĉ��c�C��9�n�-H���Tg\�Uޠ;n+<�_8V�ጋ�g ��_0���?�dvV��[�@R6.��z(�*�x�u��2�`����_ӆZ��o���;�J�gb�A�*����y�w�gu��n�}�.s����[��T�.�җm�Ջm�/f�'�ʑ�D#������>DD
.��X�K*�H��g�b��bl��1#I���R�0S�O\^s�eH�~SSSƸc^��^��8W�Ԅq�y'E$o�Hi;�/J�y}}H-O�d���Y����8JuIls��� �f������������}#���E��6�����D�����K������2V�dj����{~�>���_(�kJsraiE�rkeu�O����%��L%�:�H�5�j �O�y�������ru���q���p�.I��I5ndl,ѣ8���0�ή�f5D~G�x��6\,��3�ƏXk5q�m���an|qS��z;�2V�è�u�c�D�)�Ü����8�:K��[!?vg� ����\�ę�P3X������@�q��<�˨=^ ��I�;ɔZ��W=�⮆v�ƚ���{M9�O�~ ����N�x�.���$Dp�A:��#1[=���8����Y̾O���
�\I`�g�D_@�WLb��8����/�&WK[{���46��Џ�]^tz'P��L�K�]�T�C�W�3M	Z��;؂�&?�����4���+\������r^ԟ̛�tY\R^ �"��d|w������ơ�{_F5iuz���E���'�\�n2�8�"������ �b��<�\/�����j=�a=��XLb�^d�-fs}ƺ��$�a}z���Q�[ǟ�V�jx�E$�s[�Bd;�����I�REւ����d�������� �ݺ:vN[�oo�Pd���)�������XP�u��ˌ����D���7�����|��öm�d� -vB4K�d�X�����w%�7_�vK��|��Wg.JV��K�r�0�,..J �K<�j�JIި��>񓓁�"t�/�UD�ڢ�4�q���N�tU ��t��}�O2*��#b�8A'�� ��g�poWw���~%�@��k$�B�ڣVu+�{}|�!N���{a}����������ܚf�d����K���z{���#�S�^/��.�	r���Q����?H�� 
�
k�4+V��]��R�]!k�w��������>�n�x���
��R�q����^��L������[���F���c]Y�H���͗#�#��� 9@=W�K-����?�J���:c� �햞��K��4�����li��q��D�̸�f�C�ALTԘ��s`�G�#`BF��;���{ʼ�{�+ ���]�1l�����А�m��B⻂Or��$���k�ׄ��jP�Z;$�*��������c�Tg�7�-8�{RqT�ƕ�����u���忓i�߮��BV݀$G(挞��ZP逨�-��g ��ݺg_����l2N���i�u_�T��$)f���d��ꙿ	B�R�#����^��C����Kc�_6�7Or�>�O��F�iꇄ�C�Õ�ǗS�ňDVÕ����f�	���V�\���"��L9�)�s�2d��Ц{����ԛD��~�x�|���"�n�*o ��y�GS|���w�X@��͇��vNr�7����It��8��z��U����7�u��ߡ��4}�h���ć$��������m2dҒ4�{�F��3��i�����^��WU"��(w�f�{i�D��a%�;�>��i������5��H�!�+������R J>��uq�_W!$���}�/�G���H�g�����bN��@��-��`�S��4_E6;|�(Ib\=����g�'O� y#��,O��ΑH���� z_feM;�{p�����={���0Wr�7<��A���᯸�����Ĝ�U���DU㪧����pE���Sw�Cpsr8}��(.�s�d����p�n��M��c����7)��C%�.t��{ā�p�S���G��6�)���A?*
W^���,Ǖ�����J���!�yB^����V
���;K���2|���	���>=�k��t�W���C�:�y�H[p�9�7?���=�T%�m�����2�u�K޵W;H��*���d�����[\+�Y����p��Ntv���HL�CC��Oh���_�L3�]6qq��&��ؘ���Rv�-�$9X5휧S���I �J�(O���"�Ms��ϲ��NLL�B�ny�3!�nSn����?��Y�[����� ҆�f��:�:Vc3vK���y"��=]���������x/-#V�;B~�J\����f�%AA"���A�dO�89���X'͑Qq���{�2B ��o>ѦK���YE� ��P	��ςX��E`��׳վ�\������{Z���
�WPs��!q��ﭓ�F��g�tT��q�8��塗�L��02ח��)I����P���TˬO��V�5m�]:ӕ�.�$=�?W^�B�ki!_�(�jJ�5��N]���8w�IbŊ�:0�ZDƯ�Q3s�ڂ���>z��+ql�̰QH�wVQ1����h	%��}ՎZN�����k}��2.K�Y.��k�\� L+�~WI����Yᇳ�v����u���Z��E��A���|9v�>�3��HM�KY7B�Q�����)�UjBg7}7�d�g�OC�7y>�hd�t����l��+���1^�u~S����{Sr���t�*ڹ�����-q���-D$�	��9?�Gx���\���tmIIɮ�۪��g����n������f�e-;S�{j���1[~¦j�ňЎ� �fgm'B�Ta��#�GLT�5{4߀�k�1��2_�x���lpA5�-7E��*!�5���΀��U?��ʉ�nl~2k48L�9[�N�emgM4���æ�B�>!��٢Qv�i���k����Z�-�a�tC:���@;/�C�6�"�V�5�)}sc�L}5t��G��I�������
KW�	˗#O{�N;k���S��>B/��#)�&cUyGSSSCl�;boo{�N�?C}$��H+�4�m�7�n9L�-yYÚ-1�f�5�R+���mA��=
M8�.�_e���V���N�-��{%Bo�Z���������v��`P���w��^���K=�9���6k�h\^4�>֖5��w�?;�סSb�O��o7��l!���,���J�?��Z�[��jJy�W�ݧ�l:�����x'��B���b5��b�Ē�k����A]�y�
�w�qL�N�c���(A$��}��1���hG�6�W]�z�����9J_��7q�jBޜ�@$���@h�ټm�7)�	��z:��ڔ4�q
�šU�*8\{��o��0mr�9�(ڃ���,�x7UCV�{�� 6L4ڂ�pa�ٻ����ރ�P�.�8�1�?p�\`�*��a��s���"�G�kfjۍ�e4�ߢ�;o���.�̷�^p���9���`m�w��\���|�=f�ēi�޻nE�|�G���7�?��hA���u咠���	$U�$Yݰ��$h] �e(��QNe��l ���rq��3g�>-8N&n�i,̌T#��|����1�ݘ��8���_��C� |\	�4��M�������:�X�4dܚ5�����s8��LksP�tlM���wĉ���s7�_��<�1Ϲ"Fp���xM����k)�FXe4Л��	�5��{�-_���d��ҡC��"d���8�OEaJ�27Z�<�[�I	����G�0#��oj�\��$��LOmj���v ���EL蠉V �1ڀf֬vӲH�/@����U&g�>�����So�-r_7<�P���CZV�1U`^��O��ǬL�(�.�Ro?]%H��-K:�2�/��|R-�1���<d2��v��9C@�M�>W��"��$t�M^ֆ�kE'�]�������?*Mj\���`l���(*	~l9�����gC����N"��9��jy#v���W�P�DԆ]��p�����>_��;�����$��K�	?��I�;���M��� i��=[N��])Q�� D�)o_m�=V��	HV	LJ�A�F��(-:j��__�����>�s� 3��5�Q���A�o���O�nL���Y�p��cq~�4�-�+M��}�_�Um���ܤ0!�p�HW��B]�� !\^R7~�,t��	g�y��A|�5�[��6K���dz�S��WT+n	9h��;��!�s���M{t(}�c=G�|GBx��n�h#L��J��y���|�����_������R'a��Dr����������u%Z������g��D�9*��>����0jfg*��0���:��D�J�~\�,و8���P> ��_���J�V20����+�|/�^{��9��W�����H�U+��`
�#��X��y���(�	&��Y��Y���X�Ѧ��FZ�]ǥh[�z�	��㽰�gP��@�u������?idE���L�l?=2�\� ���Kl�9�y�bo�Y�D�Dӕǩ�������X{�UG$ژ�'|6S��T�[��<+n�nS[�C�О�ґ�
t�4������k��ٝ����%�mi�?��A˫%�ꮩ��f�Ʒ6~J��5��0B���r9�S�B"A��J�eV�P˕06J�7���V�C/dO*�coq]�)�?`�?0�m���vN�sB�{�k���{5Bt��M������v��joo��AZIA�"���j��7��)� 4������QvQ���Y��=)���?Tݸ<�z���(�� ���(˟��m��� $U��s�"*� �ݪ�}	�X�$hJ�����+�'$�������vA�(;'�;��%���5z|�Y����^���nP症0�;�����B�k��_�_�L�./�ޒ�3�~��0�n���H(�r�#}.z V� FL�,�i�7�U�5W�hu��Ͻ��Rn��r��՞�ű���w��=�,L�����ڀ�J��_/u��h����8*x��9SӅv��q�@��0��_�kl,����<N(2�Wc�^x��M��Ν-->v+�iW��R�pr���Pe�B�3u�i�&��D4�f;W�	��Q����aK��&�3����Y���ꕂ/�U.#�m�z���K��u�\�ѭf�tq� v^��̀_�صN?[8=�,�p�-D� TQ�6��q�����h/a0r:�o���K:=��wޢ�@�Zbg��È�)5�o��B
L�)��O�/�sQq�۸i�Z��8%g�	�ȩ��nyY���B|g�}�ݷ�Z-4i�=��Q�$0h���ұ�h�@��Dr�۪����VWY)(m�8.�>a����{W�{\?S�"Y�`�*C���QQN�j��憒��V7�a;�A��H���,�wfm\7�e�܈c/�7��7緬���@F���\=�Rc٪t�NH�z�dk�Y�L�""�V�k�6{*�.o+��b���x�Ҹt�:���q% 膗�.��C;��i^�8	�w��GK&� Z}|F/���h3���x���k��ѕ�m�du�!���/%⸩�|�*B���(}��7�
���c���:�7�~ӣ#d��d@$=�Hr�p��Ϣ�T.&�l	 .p����Z]a/G�"}�}�H\=���I�V�A���[vl!u���=��cQ� /n&a̶��!N^h ���2b�'��@z!�٩u��N����Hj(o!��|�@p�\�Y*:�w�s�ه�r�O5�e���Bd��֠�l� ��"��a�Mt?x�N�A�
ӎ�~R���ԑ����dK~J5fksK��3��˯ �+V�`�����S�����ϴgo"�)U���Y*�koQ���#!�$��F�O��ᓟ�\~�����ĺ����.%��%Y�O�5N`��0��r(�ң�:�&���'���y!��̠jP�1ݗW�@�B��}�Î�8N���!�_Ȑ���Y��fЗ#)�D"�I�w�O�+�P�p���F$h-�3�����O~~o-ۓ
y*��︯k�' f�������;�*���ի�k��Tm|D;_0zn�kY���d�ɬg�X)���.�=��|�K��)6�nN��֨[��U܏�nDKF���V������<��LIL���~��~-�UK�p�+���5r��F���m�?��r���>��	>[�|H-��M���[��Tw�[9����_���c���]bnY99ޏ�+^��:��+� �	^�yx]�9Lg�s+��>i蚏��ރ��M/��kõ�m��v�P���|���%S���O�8���� ��tyOKIs/����5���'"5������A�8>�'�"c��y���Hcu��6]'�&*����-�}/8=���~��=�a��G>�!���x��+��p1\=K�,vZLH�
˵i�ʙ'U!W4(��wRpP%�A]uֈ﬏U�	k�3Ȧ��G��L�Χ��oAt�TH��}�-��}�k�jt�æ������BDdP��ƶ`8���V	Ll0|٬pc)��0@t�h6� 8׽G��#mJ|{Vf���r�o�J�OB*v�<|t-(+`��0�aY�W�=�-����4����Roo��X'�AZ?j���m�2�M�J��h�m|��3Я7�8���(q�YH����]У|7µ<ΥR�-�~n�[[k<V��^�^�n�d�<��M�=��� �5�l�G'��üp0���ؐ�f�U��Y���R�=�U�Y�R�K��Xu�����b��Ǜ1���T�\}�����g�t�9rO!�#��O�Hw������Gq< �o�B� �������L�Ma��*��ϥVE��l�U�#���Q?��Ԓy$�����Yy=�S�	�kS������ޒ1�f,�R���a�S�}�~Z��A�F��O #� "���
g�V�`J�_�sBv�m�pVk��DZN�ɑ�sb�G��j�_ꓞ��ў�]Z���Hη��!��%eA�����!�Ç:c���2�u#\�Y'PpҘ��=r0��������;��.�z[lK�i�bL<P�5+�H�7W��gTU�)J~"$�6��L��p~v�~�mD�FDI���ް~�^�m��� ͱ|����T�U��QJb���Y@��tް��)�;CQ ^�k<��w��Q*���!'�%��;�"$����Βۛku[�����\�#.n�dɪ�'(ّ� �yp�}��Q0����A)n���O����I�`7' ^���>S �~�qj;�~Nb�\�?��&��S,,���M6��[�KSQ��23�2�jD_��̙IEٴ"�)�Ԝ�"�,]YHXQ�oZ��t-Y-h��F_���@�U���Q1���}���[QA���=�s�=���9o��D,���v6�w�-4	���s�$��;�ޕ;&xdR�����ba0�lw�:X� �X06�ֲ�g��~-k���=�3�4��יć@�35�^�{2`�xU�� ����W(e$��!^N������OGg�)���Th��-e�A�������N��d{<c���2���mͽos����C*�	�����c}��J���a��b�W�V��~8�Ds��f���@3NݺX
�-+]��v�u���t4Lf�M�q�����+�ذ�a�_���������%T�����N�[�:3�A��p�3���)
Mk&ثA�����ъ���l\j�� &�J�s���UhG+��3x���Go�.7T9U��|:[�����`����DJ	Vg� t��5�ܣ�)E���KI��Qk���D�
�%��q+֠!���ؒ��z���������q�Z����̭s�5Ҫϙ&|Gøn3dE�d�򉼩j���lyzd�8�<�p����G����f߀|!~c�-L�_�-�	��0���Y��~V?���?gum�p��j��l��Ɂnb=�e2D�w�{�>"�Jm�.`'p `��]�1�3>��B��2e���C��
�[ <�(���[��&�yf[K=a ��)ĵ����XD�b����n�{�*/ivB^-o�p�znGx�n���(��� ����Jct�������J�<����pÖ� pPS�q����(�3�ʴ]��<� �4r�Q���+��9t�Q��Z*а(�ji��x
<��� �P[na����N��n��x�/Ù_�Y��mj_֡^�=L�"�:�=*-}0ѶE�A�5���v6d�@Q@�iE|x�:�b����G��jJ�&uF]����Â\m�h�#��n=�G�H­E53E�Xk"lN	M��_�n�;�ZD��9߾J�->�OX��w���e�yW����'�D�V-_�b��PK   :Y	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   :Yԯ�|�] n� /   images/a794cf5c-4b1a-47ff-be53-d48f5d14bb41.pngLZP\K��%������%�����k��!����`�w_�����SEQ�5wf�����s7\YQ
��+iqU�%�W�(H�o�-$���\De�Q������(��C�����J]�%������������'www6+{Sc�Ol�ǂ�00T02��=2�==�>-�>�׍�՞��xg2��,�U<�W�"@���^����5!�%�;�nr��<넨�n��~�]z���!��ݓ
$r�W����R��Fޥ�X�C���
6}��t=!d�4�@r�7�-#���!������>ta0��ü[��'8Xi]yr��k�­�ތ�����L����c|�����ӟ�t������� <��!������J�}_�{��=�����Ds�c�����_ü��,5���kL"c��m������#o��mU��σgR$�� ,��f�h���a_a���;�х�2!�b��p<��jl���.E;�����ti���j9�_�]�'^1+Æ��ȪK��m%M��#��1��b����*���H�RL�=YөWz�\�\
T�n���� ���nǞ�����K��Z9�	T˛���2qXWŃ���p�e�T�f.5*�h��=�cPA��Ҿo�N�B�"A3�L�5�߈���R���Fq��a���4�"�1R�#c�,�����W֯�ԑ�� ��Z�꾝
Ne�7�g� ��3����Pf�3��Q%���a]�_b5(7��1���J�č`�^#���\1�|�d�^��Ex>h ���b0���G� �,=u%�
���/���q��-{�jt�l��G���S��X�f�L�'�>���Њȧ���$2!�~=[�)��ߓ%���/$6����]D���a@�U�b�1"�ŽLQ�j���#Q���х�6q)�o����&w�O���#�n�qT;*��R�����6x��0�Θ���b���J?E�d�m�Z����������]C���t���􁛢��wd���� ����ߑ<�b��J|a�RV��9u�6n��������N��tw7�^3���.��H ��_R�
b�>r'	�35h71�����]}C퀸�
�g&�'T�`|�_��9�6J�1b5�=B$��ƥ?�q7����ō5�Z�Ѯ�: ��ƬƱ�� ��m@�,���}�f1T#!�݈7zԄ*$T�� �˂��]R�H�T�e�D��B�	�G��'�^Ef����4�p��`N�����d��+p�{�t����L�ol�9.tqU�f�'�8>%���Dp��u�%]��B�0��ؽ�<E�D������M~��W��v�����L�����?PK�V�<�b]햫������Y���,^"��a���J���,��+�5V]|U@�3 �=?��M��#\��ʿ�VcJ��m�}*�x1^��O�V��Dܭ���y]���2m~�FՏ����f�8GԨK�Ƭ�eM.
ZxH�4L�a�
���t����G'�r)�οTl�U�l�/:ט��J��N`^Ŋ�q�f�$F�_X�$PX�h��n�W���ư��0��ߍ�F���?̰�5ʩ=}v[y|D�������r��oa�j/Q�Ɋt_X�mݦ���+?����x^�f��Rl���`u CZ�cl���n�{C*���8.�U���h�זP�@�2���?�2�Xg�/&4��9����Z��P��B9��˭���� <F�,~��Ұ�a`]BVݎH�;��cR��;oϔ<I���;�FY�:���!�{���Z����UF�C�:��n`*�癮��e�0\���Ԑ��\ �97��g�6�V����vs-CV�G����1W�i�)���ݶ��ܤ"���������onޖ2���p~
e ��S��������΄���X�D�p�+d�Bc���(Gc��B�b#��+��Z���F��a��T�ɡa�a~a�nʩ����͡��z�/l?d7t�4x�4t7�`D�7�^26���l*j3Lu�k*�]����43N�g<���In�|�^����=�	��.2��^½/"��\����&Gl����ܸi$wʿ!d�V|�6؈WB�a?��<����z�]�TfÎ���D��� `����a��7�!^V�e�C�_����'�`H��1�P(.)� ��T�=h��E���Vl���P���	 ���T�t�7�Tg��>G���P��ӉW!̸ �V�u�Pny%�� �w���µ�C!i��>������UV��󡟥��c�U�������J=���:��uԅ	B��ΰ��&���A�g>DŌ��:�.?�0;e@�\���Qd���d$d>b�.�39_��mqe�8n��"�n��?�?�檿�d�c�ۭ�)t�~���M�*_~���w©�{��M��pq]79��b8̕I���<d�; �ĚY}��M���֍qگ��4�r�R�о���-	}3�_j�GTP���^/��`��51wЯ��D��<��M�����hc�e&���2d	+�3j#C���!hS||����$I5T[�R�)����(���Q��."���|�B`W��;��1�z�dτ��c�|��{Z��2�CȞ˵թ��X����>���"uS��}'�4|(�ٿ?F�1|U���Qe5!�W��o:-�4[^�/��M�]����'O��\l:tR�cD_���"�X��I�@ޓM�a/��QX�"������m��f�;:�uz�3�b&��mEs����L��Q��6�~���Z��u����NЁ�qY�lU }ҷ�U�3Zhr�MP���~cK��L\ݐ���,��K�U�<�H�vM�t11�?9a
�]=�[�T�W#&u �i3�	���5[��U�dPPj급�?�B�/��T7��3EA��F�~�K�S&�S�<q�~��f԰U���[�bF���k�C����k�[>�пI�0nwS&O԰]oS�[S�L�j2�Ě� tޡ�p��Z)QRWVq���!0#:g��f8Tujʈv	�M͝�~�;[���C���/���f�ɷ�;��������K�!��
JC��(a���,hk��e��@'5�DK�LƲ��Q}&)�9�e��/����oOU����0�r-���=Rй�{3���lp��_D��a1�5��5��P~�a��j��[�,*����K(��u�i��
�>\f�X]IA�v/b_t���g=d�k3��܇�ý�	!s��
���������5|�T]m��������i�$�_c@��6�@D��R`���X"s1��X���HzL�gES�����3�7������I���g���WV�'�����&�	T3�6;ղ7S;Sf.j����3��U�T�/j$�Ai�]�1T�ru��6�ʹ��7�|��q��������ͩ_1F��枉�����](9�E�K��-遹e��*����8��.F����!�g�Cz
5q��0�mԥd4ͩ9ګI�����$�7�ep���z�F�EuY��_��i|��>H��\oI��ݚ�Ҋ�J���QОu���e�����%�/��"����zk�gT��/�w��1�Q�}�*�C����9��0��?h��-/7�:�0�~�9��m�,�W��%�"�)�I(7��2��%@/�;ʹD��m�8�j��C����M�|��`_"�u�#�����9A�-H�Ẃ�x�)L����8Q��5%(e��_��4�3ſ_�ͤ���>*�n��7X�v�����eN����nQ9����yc��u������}_�~����P�D�p��i%�Rm\V���F��.�K�c�h��ٟRB7d��\J)!a_aJ��,�&����9�}d^]\���0J���y�5r���b�|si�@�_���6,�_�T��?~��U�0����!���%Н���ԝaR�i�+r�1ڏܼ�����,��T݄�=BћOצt���!b�ʫY�@YUl��i��c�,Z�/��;�/�p��Y���^�Q}ZR]1)1����cG���/:s|.ӱ�޿b�����Zo����X�.(3�1�$�m�d�߄�?��yf�Kc@�,�����#�._�e�p����]�~�E���/qT�����n��ps�z���O|ۛ;�Oԅ�H��Oꠘ�d}��rh*�8���f)�U��Gjs^z^.#@�&��[�^�/՝�ɣ�r�}�Z[`������$^��3N�I�]��2&��3��K�.J�5�󒔅0}��lSŒQp���.E�� �l���#�4fYh9g���Y�����{��o�wz��z<����eHaA3�kn�_Q����g����oV��"e���>��HjK|/�r��rv�a��z����[��5�R=o�R���:�8v��i���g�(N��!t�~Лv�\r�L{�Y:6a���x.�WU�o?�f̩I��K6���z�.K])���BO�b��:�)@�(�	l�G����5����ƣ�� D��/��AX�OW���0N&@$��*ʈ�m���$:�и���P�?"]�g��m��-w���`�=��3�����!�ԃv�Zjr ����]�S���?LȦ���3V��w;=a��ǡͥ"ϋ�����M%�ei�e�RrݺJ�Ѓ�<x���߯�|�����t�E���J��'|�>w��?7�
3��cMS�CL�LܙcgZ�B����͠�n\���tD+s�����n��``K�J�M��$�);!�z���W�5����T��/5�9`�l�]�np���5���͝��J�=�j�B:]}Zq��2����0�ʤ�=dN9(�7��SP�������X�����G^�ѥ�`0Ӷ�(�����<��7��JQ[�4R��j*��UN�⽒k��vd^3KTr%U���<���
�,�Z^	'�C�l=�礂f�h�ky�0�w�ps���2�#�a�=�z�݆]FHi��ȹ��'��bԐ�����&�C
t��[bY
�A('�U�j�+�
H�.�{�PW�`�+�Q�_%�ū�K�!�엚2]i�w��	 j�a��	0��@n�j䟏h7v�����q2��/�k��4NL~0��wBic���Rs_�0��`f���L�Q�6qF�*n�Z���
�L2ܗ�o���r���_-������ˑ3�u4r��r9b��K5W�ܕR��~$?Ek��o��+�P�:���0��0�� N���/����[;=�e[�o-����٤�g�dP�6ܽ�f��w����?)^��ta�H#����8@L�w�R����ʅ"��$�4������� S�Lb}ȏ5=����L,ս��8����1Y�6#)�|��^�_@�rVӢ�#��V���ׅQ��l����Ae̳/)�_�O���㩸�K���	yM]M�.�xX�D���T#����Q��x�����Q<�W0L&^"��ؑT2�OYs��N ���=C�<���J�c�\�箦�;2à�=L�F�����������KJ�fRB��g=��3W����3����µ��+H��v��Y�"N��W��A����U�U6j��n̍�&�: �����d�����䐊�'�a��v�چ�	�鋌$ƻ�n%r��������+5��-��[�=s�w��ۧJT��>�Sסba��o�ʁ҆t��W%Zz=�U�Yi>q�0�%qi(��� Df��]���S�O�W��H��#Oq�ۭ�d�Z��FhIS��~߻��\G	bl+�95�h'�V�� �����s�=@ѵ�x(�i���Яr�IRa�}���r"��Y����E�5	���2Z7HP�f��^���t3'4l����^o��=�	W�s��Àp��<Up$DFl����֤�j������}����CyarOqX|"�׃�!��>�ֺ�����>�r3>)A(8g��4�X�Tϕ������y��_��Y�S��(k�h�o3���������Q s�Z���_���1�`x�'{ut!����f�bʶ (o�
�c=k�:����ǂ�
v��{��SU����\Ds�v.�2.�1�V��,ϼ�,uɌ��1�����K�@�����G���U��>zwŬ��C�]�`��i'v~��,JiUᘎ>(���$O'��
�p���@+�����6�ጏ�C��O�㴡h��,}��hz�UKq�c�KJ��5(�����X�GwU-!-��7qkR�'	vhk�	n&�-R�z�7��Ǆ�<�P!��EXj|���'��*0fC�Y9���3^���%Ud�Dr2�#hv�5��0>>�����<(�V�9b�P�����]�<���g_D�;n��>�S��xy�'ʀ>p�p���˥�A)�k��B�T��7�0D�1&\��g!����$k���'r-L�����T�!h�����d	a��"Y���!�/O*�����9w���h� r[L��u[���o!���+��)�#0|�ϩ��鼶�'n
���c L�����Z��4����I�<}7�q/��xj��	�T-7��52��@��#�E�yY9x*���si&��X��]�?O�몮��^b��anX1���L��x9�k��� �Cyܷ�NѦ1Ґ�~�HOC;X��ۇ�>��+�!�%��g�5���Q?,�����0�c[���R(ɠa�Q�yc$�	���7^�>�5]+׶hv���X`0dx�b��$I�;A����v��b�,	/oؗ�o�̔3�1����V�z ����|���qMF���pו%�5���,o�.Jh�cB���C��d�+p�cgf��Ъ�a�?*��v�*�\����c���S9������E� � 1��x���M��B�4gj6 �c�V�B�+ҕ��b�}<�s��ܽ�׿"�����(�Bh�N�|��[No�2�Ob�1�Mb!T'�eJ��oU78K]���ѱ:�v���`U��X��J��������d+�`3�5Ѷ��u���<y��Vu��j:պia0�;��Gd`{2 G�d씶��O���5�Ӄ��bh����r�Z�l,;��o��l}��ȃ��SU_�PvF
x���7���>��H����㔘�B%�;
��fQ�Қ����0=CArE�R?�A
nX�Rl��'o������s���8��:�*>�z�"���D���zr����"�u���)x��:�v)�1����TAr�[Cb%��j�J�7�4�h�|�lmME�-�EI�NW�z���Cb
>�=?�f�I���N���?��ɏU'�_���ݐ���c������G��*�2������M�P*X&�x�d��*�D��5y�04� ��K�(��FJ@���1;�ޥ��A��4���i�,M�4hЬ�>]�L��N����3�0���~
�4yWz[[[���7v��E
�Y�c*���AL�&�V�������x��Y�RKm�5�Q�(]� �n�z+�Դ؜[x��vn�W�12V���"��/���h:�Y��q�V^��Y�sl[۰F��f^��P���r
iPlk(�[����a�)�s�_��F�8�6R6~�up�BgDǗ)���%��!�*�n��i.0�^e��v{��P��|E��t����'A����j��Ϩ�:5�G�qb�*&N>�e(�B��q����$���xvހ��3�tR�n��[�f�&���Rf��No�eP�GJ�wT���'0�����.e/�`uF�!���Jf]��|�!�`0���bC��]�H�6|f@s����:��"�j�s�p�{�'<){k�=�L���˘�9�3�"-��L�\�TaB�ʰr$j�~���h������Ӹb���s���Yښg����juO�`��A�R,��� #�^h���o�~����GG�Q-f���+(���J�ASmw٢�J{	F��j�����w���U�c�X��9 �u�IV&<��y�P�\ٛ���S�FՍݹ�ػ�VB�c��ɮ̧�-�޵�$@�:b̽�ˉ�83>����f8��ѩ�}
���8�Y�ʋ��,7����"��񡵼/�K|c0,��{������H�'����l��Vne�0��?!�TN�?�_o�=6Y@4��ZyU��U��h�K����8���y��["�"�|��[i>�P��_����&��m�����,%���8YArr����x�_� ��i����$�����7?Ǫ ?R���,Wv��s�-	�r���B�YL�|D���1@�G�iu�|���n#�)[�_�(��,�'�?Yco�k07���0���h�'~:D}�d�;�]�&�f\�w�QQ�W��d����Z�rr�����~��~��l���p�铀JO��ھo~͎x	�h��`t7�uĻ&/Y��-қ�J#FY�p�?Q7�}R�>c��"�݁G2B��4�
D����;	cy�z�������W>
��&Ϊ�{��m�4�$����������N��-�+lf��Zw��܄� �+�@�ݔ�2�2T�t��	��h��O��*��!|��팟����L���)h�}N�`<k>��e
�����pu��'Y*:Hy�}�	���..�fu�E2)�$vN���Կ!><��)�1{��"C���u��Qc���+k%Q�Lزu�p�ML�$HDN#Ku�f5����(��Oz�iT��H��	WO�V%��j<R-(����Y��a��ȉ�x(r�!hq�[��O+.7����5�9�A9N�E�}���H���C������$��5Uj$�Z�>��Dbv=0��u0%B����cm��t}ify8O�c�Ds���闶e��ő�E+��w�2���⩈�z�z�;�ր�:���(��itDO]q��_������PM �#k���_oư;E�)��)��X�����L�2p���j�EVw���#ȸ�=��xH�rQ�~�:��Y	6 	DaXP�ච����$$*�dp��~������J��-ʷ���:��}6�cJH��xw��̌"�P��De����*b�d�;���W.�6�i�~��C/�\qFe�V��]0zby��16��3G�z/"���C?�A�	c���b}�'L���,d��Ď7L�l��3g�|�$-��_3�������yTSJ��aw��ƏT� |/=Pd$��V&��mZ[O/u��^w��=N�3�KZ4n����C�P��9�tC�`�1�5��!�lx�w6=��c7��{X�4U4/n�>|��fY�HH�lz��i�3��3o�@��v?d�<J��j¦9�KRu�wRj��v:�b���Q�^�`�j��$W.�0����	�o�Z�k$A�����ʄ�:�ĒF!c�ý�i�h���`s�y1S�_^��"��
5�
�
`�{	��L���ch)��G�n�Ր����~�[��U���9�Z��;OD�jA��,���K7�铨������"DL�0�7�u�����oEk�\�5{����ޫ]UH��w+N��Ӎf&l�`V�y��*�<L�]��n��h��#j������XR�u���Ʃ�۱RЁ�@ɟh�
��E �[@k��o7;���e�R�`'���R�Y�9�X	�nƙ��,�K<b�r]�<N�H�����CٙfC%�v6��.8�ƉEb-~�*Mih9�H�J��������e�O������'T��� �������,F�x���6��O��w�5�;��vhzY�X�L�C;���v��9������.���1��o���p��0VN�9���)f���BM��,�2z��3���Eo��R�J��ߢu�l��;J�p:U�*�Z��9���Q!�e�V4��8�����[���Z��$��?���M��y��'ؘ���Q�>�L��4ś�U!JL����u�$�>&��=F����}X�""EN����XɸŢ/�7K��0��Dq��S�ovmP��Ab�J���w�~J���8cÉ-?�#4;���[�A�-���E鲨�J�_�bp�w����p����O���'��Z.�T�a����ȁF%������*�ሃ�#DDFŰ�uuf�yff�'ߴ��7��2j��Z��ea$08�T'L�������G�M'�Tq���p�<_���D���\t�l���U�(a�ݘ9=�?��Vҫ��z���Z��ovvïP�wCJD-O`�;�XC��O��T;k8���`,�w���d`�`�~��]�r��O/f;
x��v��7Ӝ-�b��
�yNMz^��/����茷o��",�\(p
Ii�N,��_�F	]/C�̩�Ւ���2�H�>�u(��6\��neF"}���@IO�wCP之!w�_��^]i<�cŷ1���C�yG
�%�
ߗ��jH�����{�#Bpw��Ҟe�k�j�*��\|sKw�u�,��O���<4���V���V���7�{#�V>��D�I�����T��:V揝J�ku)�Fځ�:�ɇ���H
}nA��vxU\��boo���^FH��5>�A��V�_�f��
_�g<8x�Uax��	��|֢�N?x�d�!��Ԍ٩�6��_�v7�*��XH�qh�����v6u����L>� z���q����\���U}u@��f>;{S�	�+����q�&�JY�&��_a����<uY�@�f>ݪ|ek'Se�B�6������ װ��\~�P�^/I��l��|�ǳhsh @{hC5���Ϻ��p��$��p�����K�g�O�4ve#����vk�P�����i>��ƫ����躉��Y1���_���zde����
,#s�qc|Qih�U��)��˿Y�iyl5�3C\����ƙh��c�k�̪�Jc�7�����^ONxl�����ܡU@ȟ�ށ,,��IM��@����j3F� �m���΃�g�
�'�M$�B�V�F��N�G_`0�?q�^��/l��z��4ts�_��o{�~��ѯ�=�e�'7��x~��OWR��tP�BP�8�����T���9�@��v�U�!��}K��;���Sgg�ⷁ�r�du�a���\f��R��T��]�a]��m(4��.9���pX���WEpp�f�����mO�� ��1��;I	s^�a��L�s
*>�m�LY��y6|sI����q�U�|�Ri�뙉K��s�yT���r���	�X1?XB�cpxU�r*j�bT��BR[M8�k�;j�F��ɀ�9�pȭ�bAO{��7¥@,X�է���.���q�TZ�V;������!��(6І\���6�f��ß�!����F����Za�3�+���}��#<w#h#%�M�3�~�l�x���v��uS:&�ue�W&V�ҩ�<��(�n���m�bwG��ʆ�����9�pGݐ!;r��a`}�q�ي��˂�T����߮Sn�eA��JD>wg�������^!���Ԗ��ē�V�D�U�}�!�z���j>h��~��ci�}�i������揞
h>Vfd�>���y-P��A�0��&��Я5=��jU���)����B3��j��W�\�E���Y�兀�Tx�v�3�-Kz_$wͧs7iy�SS��>���)ci෬ˁ3{����Ó'ӡ'��ls���x��1ş6V�g~ctP0��ɡMV"�3�)F�/��pv��/%<ȧ>��p�j}�Qq}��yL�>��p�s����R���`��w��M��� ol���B��c��N�I���z}<�e�ل '���:n(��}';#��|۱=��bm�� ���s���ܞ�݀
O����r �ղ��������k�E�3���Њ���\گ�<��<u�h�;k�u��|e�|�B����љgHy�����4����+p)C�J��6G��|::�W���˞m����Ku� 
H����>�i� !QK�O�o̊5k��Ai��sy�M�{
#��9��E�� �� sB��dh�����9��^wT����)�C�}8���,?o�G��Iι�1A�6v3�}�t�ř�"|�M
i��%�e���e_i�H#+�Zr,8��谇�{����aiLn�0=����}|*��g��1�͗[.s���D�8�Y�Z���.�a�O�ƪ���%0Rj�#�+��|��{0P�y�#�v��<������.���P_����][�i����U�" F9����Sɝ������W�@���s��f5g�/)Ik-q汫WlZux8�Xe+ �3�,�N�}���8�:��]7�^���������rz���U��ߏ�$��y8�@�:�ޟ;N%Fn'C�,�=�U�,�jW�����9�����b���p�/�'Z�Omt���ھi+�Iqׂ�Qs����k7��.A%�t���|:Q���V��.������Bm�l��|�tz������^��KaRP��|���ERO�����q���w�XT�n_��n<�5�9b�9\x����{rZj����
ce��zѕ�`��5�W�"k*K(����|�wJxDy�<|����rr�G�c�6��w+�q4�O{K2��d��2ZY�*��Y���i(���\����ZZ��e�D�3�%R}�7����,�g���+C�EL�.��Y�3*��g���-��d9޷Ϥ3:Lo�g���U'|�G��f��������r�9QDD��`S��9uM�p$��$];��?2C4��Ŧ�VI���E���
Fi��~�G�g�����h�-���XK��c�}&�X��}�a��g�)#��]����p0
�����Z�$[;���+t�O�G�JM邫�.�j��	��16��#�v\�X�:+�D�<���~Jy���R\��?@nC����kJP��n�+q��v�{Yc�ֱ�d󂜈x�����yi���8I�K��]�W���)�w%'��p��m?������K"Hc��ylJ����۴�)�Q�n��Ox?bǜ��7��9�mz�f8pE�ܽ��-��wS|B��Qs�S5�+�^<�0>[l�#$<T>~�;���y��|�!���J${�GM$�Û�M��k�'s�3+x�M�9��$�v��ޱ��%���>_����:��ޡ���kI*kM@�^�q|�ỉ/1m��I[��l�%�O�#q���1v�`�]��!ge�`7�K.j�>��8�CR��l���'�vɖT�������A��ŻP��A�Y�)w+��~��Z����C�C��>y$��a;�be�$���i旭q7��Ճ67��F~�Uw��p""O�V��4~��%��.�i��s�}����E���R`d���poU��* h�V��f b��q��9�MM���mJ��C�O�|m�&5�<�,l�̰��
� �]^������� �H�z�"+Ҩ/Ι=���I���0�FکU7
����bְYu��p�ׅ���P�e��A�iy�?�u�~��"�N~g�輝����і^�9ʹ?�*I"��P#�3��g<�J���f�~��Ƞ�>�q=���k�Y���,�~l���"��ԩ��Q���T�W����.�RR���;B�����M�U��m����� {}��a�7)r��uM�zVHT��d�w��K��c^�m�C�2y����8��G��R�h��@GW��9{~!'���@"�=$VzA���&�\�
j<�����`��K��],�5Q����4��)����� ���Ӑ7�t#I ����!��[`�s�?#&o�]Vo������ư��XqX;� �*�gTЙ�l�~�7^6�<Ӱ����ۛ?���&Ě/ "����cos,�E��'�����h_9�<�*���x ��C�c���M���8maWeC�a�S��UI��+�JS������䭝_r(^3�#��t��I�>4�p�c-��"��F��bb���ເ}�Jx�O��0�7��<�g=�o�P����S�ԔX�}�������q����F�Ҷ��:D�z�$��w�T�����)4�����.3������D�3�L�g�J����`�#�g�����;�P����@����J�.��-Z|��c:��Z��~5;�a2�V��$��rd����T���Y�5V���cJ>Yq��T i�Q��hhT7���YF�2�z�MOOX��W�����e�iy0�Q��^��^Yvnuh�C����r��uL�7� ?�;U@��B��N�Ov@*G�l�L�KZ븖֙s�9~7�b��#4]eJ<e-G�c�Ƞ��ej�͡��!�~�}���N�o���f�"P�w��Ӡ�]Z⣗d2q��n!��4���ھkOws	��xj�wi&�]}Y��l6��'[�_xu��5�y�'��V��l��cO��P�0��y깟�Ύ0�~L��8W�{�w�3��Ei��&��B�Ʒ�w�&%�z�`�����t􆽤W�-�ݮB���Ba������Fqћ���)��bB�hhY�m�^��|s�����nH��eX����n��`��t���ؕ,OD1i�.����o�$[��9�p���x�ڨz���Uo�^v��0muF)�H�A��:NG?��n���xu��jG�l�ق�~I4$�P�����c�۶�>����}��$����qj=�ܵC�ׯEwЎb��M4�z;��`	��;�"����A�x�F��v)��,@em���b%��bk32��fR�3�y/=�q�t�2�0�'���D���<zV�B����c�q�b�MD(k���UoUag�c��a���R�͞S�J�����ޭ��4W8R����.y)�r7A{�TC?m���LrkU%��Vdg�<��	�Vx��>~_�j�y�H
��}�x�MHi��f[Q��6(��:Կ 5�b��C�;�����0���<��G.���Q>;(����2.O�y��"�f8�{)9��G���;<6B��u�U������y��D�@�LΞN՜dG�K�lh��m��J�7W���8��!.���V�&��'h��L�y��g��ޯ�r�юȰ�{���ͅ�����캩�p�dl��
!N�{Z�Ny��i���L������c�U�6?9��aL�7��$��X��"�W]*���PI���PcL���XV�9�n3 ����F�w���6τ3:Qf��O�(�Ԗ�~�z�7)'�����|~#����H������Z�����/w�w�.ʐ��A.c,�Y���'..Y)+sP��^��	�?BKCw�3�gu�Ʌ PM�O;����ص6w�|ޝ�*_ʈVKc��#WeyiHqg�i�굝��޴A1o�8��l�k��!�<�m��(����ruQ�h-��_�S�?�a܈��v��e&�wp91�C�B�K�׮��#5v�Nk6�t�G�hY,����ϵ'�`�۠, ��NiH�"l����ڄ�i2Կ�_�J9: ĠA�z�P�lTん��ܜ��=����N(�$;��̇|�����ݭ���q�UYh��n�{p�I _���巀(���8y�{�_5���̞l-�t�/�<31У�*j�?��Ch�0�/xr %MOhQ�n�ש���.\@��a�e��y؉y�kg󃵥�{mX�R�h=��vJ?��.X^{���xRQ\qC����1m����U�%=�����{�7n�h�bm��;��Nt�h80������eL
�|`�5�~:ҡ�R�ٵ(������S~��Ms�9
���2Ay�|��ԙ�P!�=������5}�4��msl�h�~��ja[4ͶlW�$�.�����J�̎Y]�x��D��^$IfD��'x��xp�Hͧ/l��ӽ�y�|����N�s�J�K�2�./O�;o��.�j��n��
�̓���r�B:/AYMq̻	Y���Os/#:��6d���;,�u����[���/���a�y7@��)���o:j�����yU��/j�R����1:[��;�1�~�Bz�m���wT�|�8��]*k\�n�n��wI�H����ٶ��-}�
O*n�#O(�_PB��":b��8#YGvlv�%ptk�%�Q%d�&�%������؞���IK�w��f�$˲�0�/TN^��۬���g����T��nD9	<=2�ޭ{����~B���o�6��k�V� ;	"��JH���0X[�]�
H>v艭Uʾ����[�u��:a]A��jx��}�\h��+m�����>f3n��;�5���S��o~q�)i?=>�d�d��7l(,}�x�-
�4G:���<YZ�}���V���	�LP����6KF_���ɮ3��;�4���K�E������$���GP��4�;������^+��/�嵓�J�s݅���=�"�����ō���^)�{;X�%��A����]�F1�{�=�wt�!���͜�B�<�_�T<tg>Y��@���.0����u�|���o�3m�	�~�rIf��!�i�%rW�M��ə�3	}��=���L�Q��;y�螒���e�kJ��Ի���M���F�Sa��C������/@�9<��ܣ��O>5�U�a�Y�7Z�U��Z�9G4-�4]�I���M�#+(w�z'�_	��E�����`�sy;��If*��s�����1��l�_��nԮ=k��5j~jo5b�g���ڻ��Z�k��(�j� BIU�Ub�=����_��+y�<I<���9��9��ۇm�KI򣏰 ����fqu��mʍ��6�y޶��H.�.�x^���!XJ��q�I�`��KR	�#��6f�W���~���%�g~�T^���5�����I�r��oʯ������@Ȭ��Վ1�� �f�~���>�����v�e7%#E|���]�C�1*���6v�25N�œ�	X�t��5���٥a�w�>�)��pc�y,Co��J�ϡ1�����*S��;x+�L�5�����DY�ê͏��v�b��7�}�a�	�7ؚ�IK��]Jv�T���e�8w�<�8�?}]�����6�.�Ƽٰ�(}O��"YBy�i�iu��2�/��藨5��v_=�BД�S���</_���[�wgfZ����	\J��q:(���Ҕ��|���l��/���b l�v�?I��$3M���R�M�C
v�tf��� �7�Z��=(�����
�S�rY�4��p-u�RE�KIgN�dmꘜ ��t�*ԋ�"m��(������ 8;0��5���FidVXU{}oċ�Z���I�v�)]��=q���o�p�;���~�&b?.'Sq^��_X���t����׻�=��̓���r�����6.�fu<s$0�_|��usJ[xA͝4{~�pTV��c�K�M��c����u]P@����yd�(������͓Pm�6���`���ư��q�E�9H`�4�HG�|�S�P#�z�$�g�9��$~=I�k��5;����]�' ]��\$���������EAѪ�J"�3��w�n�D���7��zi�\WƎK~Ζ/�h|&�?X-@��s��s���C*n�xY��C��t�]�J��%+���'���;S3�h��ܗ����X��:��Mw�T�qz8����^?�q_�'e��(~?ظ`|����{���a�<\%�T�i�5���cv�f��	��JY*΀a�MI���v+�l~��G�^�����E�|3�/��Z���%]e|�R�}\��1������7���~��笏�� Of�m�so��	�=�+����~L��8.�߆��$�+� /¢5i�^�=�a�����	�7߿Kᕠ	��i�׸��n8���`c���;)e��}�,D�.H�%2�����&�lT�F�+V�$����1G�(��̨����w�n��q1C] ������ޠ�R�R����T���"w��e�W���<۩�"�&��0f>A������n�^N=V����j1�P \p���TQV�Чϑ֭�)�#C����=�pp-��e�M��l�G��kpz�S躩7h}��H]�%M�}<�,�^��V1���Ȧ5��Ƥc�.�G��2������,�}xk�<�����}���%A��Xf̍d�.H��W��oe�e�!�Wp���'�G����ŗ<Am�������;1�e��]�tU���L��."��Q�i����r��P�.y�j��q��x�{'جyJ�.�v�;�O���x5��@@9������kp�ZR}�"�6��Nv���������
d�?２ٸO���:�{����r�aB�^�Xu�p�yw�׫'�"�G�o����\�!��l�D�� 4�>o6�!_��P`��oN�d��n4��n8��5���!����fX0݇j��*0}O��GV�y���ZCׅ:�F�"���ƽ�Ӻ�Ͻ{�z�`�E��.̕�-7�-����7۱'��s�a"�s+�F�\��.t#�tyz�*��V�ɔj��q�-��9�C�<�X�c���+0�JG�I�Zo�ius�Q,��q��Cb=��9��r��R�;��ސ��3�N�
!ra�m- ��q@��(x5x#����{ �!��~���⫟���B����I�b��� �(E �1՗�kmJ����$�(�N0�K���\��)����W�1ڪ���N�z��/2R~v����3��Y�m����0�Ѩ�%�|���i�`'2�9�'/�?_�#�`�_��0�jD� <�'���`���zIHl�o����:��N⏂|~P�H�[�f���d[r�A!�yAx�^�'��� rRn{6��o#[e�\�g��y�1��#j�>��UyۺK���� ��=k���$��,�=�7��2���ϲt�w�a�����3�.uJk��]%Z�V����)&*fH��S�e#�~��N�x��{����x���2���8]�2DX������J�Y�27��v^Ǉ7mД�t�q�\����XO�.x�lb��X�jGyX<��a\����Z�-�i,1*מ[�_���j伂�}o&�rN_.x��l�%��kU0(��,�Iw籫���hӮ���ٌ��B�p_�hx1O9B�MX��\G�-�W���6\�,7<+��$A���&Rl�/�NPz�c�NOwR�Fϻz]n���w�h�L�MXeNe�{��%Z��䩬�S�`��h��T���T.^u�0;�?Sq�Ԣ�3VM!�{-T�{�m���Н��&�iư��R���*3�EdV�f�N?]*��x3�6]�[b�)�Y�p~�I�=4����i����|��=&�2���M)Y�$F_#{a6�@՜ �P��5��w�%�ռM%q��~�M�D�
"i#g�3�\ ���x���n�j�䴭?l����'���XJ�wamB������v�׮ ��B���BꂊD��>k�$s����o�u�+e��c&f~���Q�u���"�B/��t��j�o�@�*�5�*�c�y8|��J�iz�i�\s����7��ջ����y�7�0�Rf@�v��������}�E�F�/ۡp;k$:��F��9݄��9�/H?
���p!ҿ��C^^�f������מ�!�$*�d飷��)r��`'��亃ЊZZI��r9���GMmE������<&��㦶�8(^�o*������[�^���%9���aRL�ݓ�}��WP{q��	рR��� �H�{����q�7���E�O)�u�:8[}��x9E����k�݆�[�7���O���*ɮz��������ޕ�/�?Xg�^&��<�kUdv�9�&�>��A��l�o��V�Ud�%Q����e���E��7��S��
�Ưx���	x��<����?54����M�${K- '{����Jf��h)��ѭ����,�J42c^p;J�v��T�ҫH��]f:�������P?��
�~t��0nJ�+.��ǌ$씄��##���1�U>+c�<f�1�<�L��x�/�z�#yR 7�R���q�/eY���#���,�ٌ=�K[	��)�����}M��v��[n��1Y�L�T�.�݆�=�V�J y��)�[��1<�t ��:����8촆�o�}�p�Jΐ�6 Z������1��>C��S$7�[��2 F�� 9݇B��T�t~Zf�Ӊ�.�s�Zk��'�P��nZ���Ǿ>f���]�VLk��5���*����J�Ƨ�����}i���T`�V���?�CE����_Yi%<i�����+��k�S��u� Ծ�*X���/G[-%�Q���r%Z��ܻ/������د�8��/$���y��! j��
��m�pt�������[�Zp�K]��J��
{z{����0��q���!���m�H��Ϊ��W��\� d�]|i�3�&�Aq!�`=��f��t��a�����IEKd����7��^�${6*��`�ʹ�L������=(�-0=�#K���&����pbb"A��2��o���U���E\������^ʏ�����^��v�YHjn�A��v{�}��R��aɓ�3�o���+�偬?�q��g4b��&�{�uk F�#+���fۿ_�j`���M�	�J�Q���װZ�tS��!�/F��%��=Apl#i,~�� 3��/�=��ص�64=��2�F����ߓr���6��%�X�����c'A��1lȷ�`����J�\\\�e�=tҞR�F�(bO�������`>_.PC�����^ו�̼?t+}4Z���j/���VZ1g��D�Q�W�,�r�=&j�=�Uw��u8H�r�dڢ�G}�@��Mڨ�9_��\?�L�٢k;-�����w~�6���35��� ���z٣��H�OBlb:/��,:���,������1��b-w8*��(u�����Mw�=�v0	Ag��ފl��ʈB�lu����Q�b_����JB��\lvz����f�9c��<]�,��$~=h��SUK#wj�)�g~��W[Q�䩄D�E𞈧إ��e��Ç�^p����<��9��Ϋ;���fh�|�'a\�a(��Q�Zo[F���̦���1�8���I����?aO����1%�tXI��^\̸*TD�QS�ٵ�F��ᗃ"�,�AJ��]g���]�k��.=OU�Q�~A����k^%���������xr�)\���U��q�	S:Qj�Lݓ��J9���B�A�J�\m��
�STi����p�3 Uw�6��s��/���X�C���;8��!.�iAx���-�`�ë�hԭ;�[�,@�HPf��_����G�E��}�+o�����yU㭠_��!d�M�E���o��nC\Z�������%�OF2�%	�F�k���Nn��N٥�c��#�x�HI|�&�1]�s���b�?5+��5�2��&�QY%q<L�!R��x�c�Z]�&mC�;�Fv�k��Ҟ�v����1�8�<���T�_��T�,��nd"k���:f�2�){�]�G�������}�v�9����Ǿ�L]h �{�q�,iϣ�y�h֬<#k�� ��BB1��'V�^gƎ�]��}�����;~�pgC_�~�=�f��f1"9�]�`���v�U�7�)��|��W�N#o�����
/ ���<w�
O���!�X��ٍ)�l�b�IUr��G"$q!AB�<|�pyk��F^�k9����tw�S*���ti�Ck�(���M[i-N�#�͊��R�V�z
W�@�[k���Ϯ���o�)���4A��ߙ�WM�c(��x��Q��/�J�OK����ށ/t��1v�̈����X������j�uߵBr�?@�Bgv�*5K�d����>[��ET�[��7��XX�Ot���/$֝7�#+�Hq��D��n�:r����o���������R��ba6������΢���Vw��psy�z$�AIdā�i+���1i�8g<�����`أv��j62���s��Ĉ����c�¹X���C)&@�`d�@�)`K��!r��c5��7Ϳ{K� ��*J"U`\oD7`��Y�w���}��JH�\|�e�3������}0œ1�/�J0T n5��wBlA`�n�.!j�q��*S��z��<R����{;�ԫ�W^z�8c�G�,�b�r�#��/�	0������~�Ԉ�>��Sg᫯��.���MM���r~a��xg޴?BN��2�s�q=�lWU�0�:Ǭ�����4���'�,�~��g[U�7�g@ Cxw0 � �k�E�$�E�C-rmi���H!MnsO<�[	�nd�U,&ӕZ���C�Vқ�>1�#w�M �I��6�|���ZbQs����7��_3�z�ɱ��~�&D�Eܿ�֣�!0T]���%pG%�(��n���W�B�o�O��|��\�Z�'yb�\,Ik{ĪC9s����u9@�M�iw �@���A�;��gW�K?0o��s%�<�i�	�U���u�A���ϸ��@�@P�����!�{�#I�I=�T��8�L������y�~�o-� 6�������(���S��S�~��S�Ѥ�	6|��5WI�+{���^�9�~o�)A�<&�n~0�$�?���y�j"��_�}�����[��+P�E�ɜIS��t(>�	|����6���� ֜�y����uOX�^DS�x-��^0���a�﫻!�񄮱���}�WH�ɪ+���564�ֽ/��K5�7ԝ�4,fUW/��=����g|ĥ��L���f�<�z��6�y7C<?< �����@LQ��&�@.��魕pPC[>�,N6N[�;7{e��7K( ����o-F*n"�F��R[���∇~T6�ܮ5kQ�$�1]��2H���4���ϑt��h�
?m�������%�-�9����jf�;���74t�׷[�2�WS|+N�O�����t16����[��
�S�+'ߍ�K��{�vS�zj��!�-��1���4l�q��=��8�G��uu����B=�;5!��Xs�mEc���ƙV�!�r7��,�s���1�A��0X 1�Κ��6�e� ��Ժ��,U�p3�f����##��>k}R{�C�^�O�?<%ЭlZ{�BBqj}:��5�J-���lk#{,.���� :�B�o�(>��!	,�i=�TT6=��9�\r�py].�HJ-�Z[5���E�-�O��:?k��R-�i�H�~],<���yqf���~(��ړ��P�,��������&�����r���t��������E���a��Ѥ� jd�;������&^��`ڿ��
�8��`B�L���8<���B�]�Ģ�ҧ{�]|W���ilS]��MX[����&6�5}��zr�@�%��oX�;\UY��>��e��YT����n��tBn2W�*����P�+3 k#��*�񨪑aGɦ7l���v&���-g�?ۂ񽺪��	}E���P㩻������zg�$��\�DLW��H�z�qѰ� �=wHid���1I���_#Ij�jC!(�$��L�s�\���8��mj��˾u�*L�*
��]��Ө�RWU5�d\a�3a�Y��� �S�ț��n,���~��3g�k�6�������%%-�I��M>�!�QES� ����S>_"g�
���HO����h,�h�C���5	�gBݿ�������{C�F*t�a���N\�u��ʓP��H�ҾL��G�����λs���DB¦�կ6L�:�`�KE�h����hj���`����W`�%�<���(9�L�~�=3���C�Q�� ~S�)��ǂ��񐭂�y
���ݫY�����l���@�v��h>w�#1��?��j�:�u��ެ�p� ���<|�'X�a(�1<7����S��j�i�;Պ�d(�:������6�LP��}�פ�ִ�3��r�6����K#��l�&��}����SO0?�،�֖!8�r��p������m #��3��r�ݗ�',sq���/��TIQ��O�S{��G�4~S��|$�%�fr����@��A�nf�n�����xmvG����!�Õ�)�j[��<�v0�aPtq�NY��X B����)�F�o�w��/0����fr��\hx��F�q��kl<l���{n\ap�#�\�#4=�,�w�+��4�
��Y�+j��?��6N�E�̀�	�X_��Qw2�s�R�v.�Y��7}�0p��Ƨ�����t�P�msYId�f�l���������U"�=�l�����g�	��n�k�����a�z�c�O�L5Ds� *�(6)u'�>�`�����n�4]~�*[�9-G�~P��S�؀��tHn�o��K�N���B�� �)�R;�q���[�'o�>�-Zf���j��/��[���X"N�ח�y�,]P�$x�b���
��(��כ�5�%݌��?��P�~�����D��'i¥����T!^�:����,U����H*e"�ω7�w웅
���S8���"1��*>�>H<A������/��<���n9���ż�kj"^����}�D���j��9��㭆29b}{�;>�elc
]�L0�P��} ��FR�)��Cv�pg���U���"������>�H�hT:�i<�n�wŝ� �o�h��e6F�|h���55oк}7l���?b��Iv������j�bɅ�h��l��n�Ϸ�y\����^�RFLXz���> $~VHc�{�R����H���@�Hm�5�4š##��f�w+��f��������94�nh	td�b�U
�a�8�S)��|�0�3�$����Wcڜ߼�2ߟp��#���&�J|���(j#V��N�]
D���4l��yTs���Q[�a��~�p���}L��'M�����k5��;� �h}|{p��M��(P��c�I�kA��Q4�!� SNSx�����Oڇ�MW��F��m�l�\E�_���&��|~�K��5'���E� ��˫M`G����*����%z�q�|Q=��f���<{������K�h�����84�^�L����h��-�q!ʇ`�N�>��^�v:�\2L�����7:�8���Q�ؐa
p��0�J4W�O"��bW\l:��������3�t����}��;�"�E�]��"H��ocV�˛���g��o�����8\ԋ�Ȧ��	F=Z��о��ZRn�Sk�t�9	�t�TL�<	���e/�Pd�>&Lj+�0������F Y�}��/�J>vu��~�~suus�az�b��|�U^^X�/gP��^��ay5/E���Y�xqU�FpQ�?����>�=t���ܓһ�Y��ر�ȝt��3�����W�r0���s�&B2֣�x�F�mb�k�Y�5o#�TD�gDuk��_'[b#`�0��}gӠ"\�ۿEӁ5�˳�{���u����Ӓy�"�\��>}gO{S�d��ӛB����^��[Z_?�n,ˬ&�_����SU��J��m��h�S��G1�,J�c~���;]�w\Y��}}���%�ŋ���TBK�x�x�^���yM��r�:@0G��K��+�X�C�p��m��H���t���>�!b��v��}�2�-(i��l���"
\d8G�ÙIO�92�?�LI��9���{#>#��[ؙC�Wz�ѯ���k��r�- x����◸�����������q�=�A�"?��S��`T����{1�X��&��������֮���{�@(���Hx�$�A� L*QI�ݩ���}a�v�N�EZ+ԋ�7<�.LP�BV���cql"n�Z[�\v� �7�i�>p���y��v�������6=>��%fGn�K�2�.[����>{b��\MD����G%�h�'J��#8L���=W�+|��X����mt�`ʴMԪ���;MZ8�� �ŝ��W���t�ᓛ�������:����R�X����M�Tǒ����z�F �c.��`V�FO��Ck�.��{7���w(�3���a�}�4�B5E�n5�a�z�Xe5u��EԬ�VR7��Z��G�F3�rp�_�����N�@�{��6�O�f����[���S�H��T�RX�sqz;��D	V܉��mi, g	�����\�߮R������E���wz.�H���N���������y2?�9b7��(u�1�_�KM號=M0�a�~�8���0'��3��xT]���$�\�^��<�($�͙�5kx0wm�ɾ���*�<Hޡ�����w����C�p�cyd"+�pgj?{J���e��wU��'�)�(��
G^��*�9)2�bH�]���7�@��4�bc��B!OST=��$X� �f�G۶�1��l�X"O�#N�\Dw������P����!
%��A��'yF*HТ֖ �[x��`|�<�2�B*0�lk�)�7�ʪ���-��&� fx��@_l!O��`��a�0�+���{X$μ<�,�;}@��(T�JF�YI
���u��Z��759�^HF��Qˀa��i����{�㠸XG����\�'wr��-Dp�+����0���,�pn�q��V�B�l�^Qv�^�]eh�r;|R嶠�X����ݦ���k�"9��E��[�q��-Pꩇ��h-���rZ�&Qv��y�k��	��Orl!V9j8H�/�6��{��3wO3�M���wK��D�Y���O�;o)\��.:����D5�4S<{;�y�h�Zg;߽a�O)�H�pPt�y�4�Y�wf%�bȓ�7+�Y_��#�m��QW��B��BM���nkdj�"̊�b���qS[br�)�CA#�Eb�D;��C#ܶqM�����)9�Ѵa9�Rͪƌc��H��_q^���܃�'8f��yv�.�D����H1��M){�dwz|���;����zC�K����,�V�TB�ar.��	�%Mm���[����@ZqwJ��K����y����A�d��/@�����T�������`X���PWF1'K_]��;�����V1q.AѮ��+�b+�`+�������ѱ:���M��A!" vყ�}F���"������%�AL��[���sU�FdW˖���[��|jjj	~Ƹ� l�x4��r5$n��;�U]n�l���v�.�V�uِ�$�{�f�0��	��g�'r��e0S��KFEy�*Bimuu+�O��A"λ^q�l��D}�gW~[�w �؍� �P��M�/5;�u"$Q���<L�T~J�N�$oo�#�O�����b���Cb�`5 �SH��:<�m�vJu(�ڞ��Gu��ߔ�4r�ݺN�&Zm��̌ � ����,���ț�X�������?+������P*�@��t�]�G��i�m
L�v�׿�d�/c��P����������w��&K
�f~������
�k6���������󑂷P�BW���G�t�,E?ah�"++����Z��0� ����P���v)�k�Oc2�ޤX�Rp��%���w��eq���0�3x�xD�x���%��J�u2���O�����������u���b��9�r��L��O_v;R��Q���&�oi4oA�zu�~}�����݄����^��4x��l{.}��1�䫎��5
�����0���FCi�;���D��
~x^i��O.琛+�����I=�+pe�<�i��=����a� xq�1���.�0R��i��_��
�v ���u���7�!`mn�i������������k���`�\x���|ӈ	|m��K�����vr )��J���M�Tg�L�	��M�*�n/����.����k���G���լ�X"nM�X����pG��O}�$:!�R��\4F�)�y^\�o�Ro�aDa�p��D�&��R�l����$kkj�\KgO()���#�����W�=�'�c.�<���t	ɷ����i�Un�SC1�����`�ռ�\f(��������&��]��5�oA�y]*o��.{�� M�I���~SjR��C6��B45,y���k�P[����+�qlCp��fOq�}�*yR�l�%�̺8��şNrP��*>�f��+�ٕ�:�d��9��/?�|��d�#C�ߴ�i��2C��v7��Rq�����#7��8̘���c� �p�eI�[�N\��~�w�Oo�}���Wn -d7� 4)���[�Nl,:�V�Nb�m']�[^ �4;�G\����<��{�8g��::~���tR�Y� 3��K4���d���
(�x��kg/t��pU]M�]�xQ�E��)6��z�>#N����gv�ɻKfǣ�{�5
6�+�V#�ٖ���$�㗭L����؇~�n��j̸�����mq� g�&�^��2��Cx�f��G�{�� %���%cZ.oq�)U}�83 ��R���tQ[]]����1�ȸc�҂��Á�m0�~������v�,�O����PvK���wާ����������#�5n��
7,N�Sa�\B����D};���.Y �����l��^d�ήY�\cSVC"� �S�~��'��	?��=U����O�e����s���%c��ȡ/aXrm�-g F<�n)$��p��.��$߲���@aq��|K�٭0��.ƾ�>K�1N\�����\~�`l�����4���\(�O�X|ڰ�ӑ� ��r�=�� �i����.�z���6��)���GN��/o��-�]���,�?��Ͻ4ă�
{�>�'QLy��X���Kc��-�e��sFU�t��4����{&(P�)[�KP@�v[2Ȳ�ɡ�A3�4��]�q���Ⴟξ��ʓ$}�D�����~��,��zD��j��z���ӟE���'r�0FV�'JS��G��&"�F�b�BM�ܞmF��V�c� [(�P�w�SZE�9j�,���r"IM�Go�Vt 尖���})�;����t��QEM��8�zN �ˤ�e����.b��̬� ��UΡW�����I핏Wd522�It��a�uMu��9�um<s(�7t���v����:��nꔊ@�|�2�qh�Y��L���D�OdA2��V���Rc�9",�!�R�Pį���iX`z�3���oqYC�(uf!`�)�O��j]]@pȟ'�n��%������,�Jci$��5MM#j���^#�>���eV�Q‗�h��y���HL��FY"՘_r���] ��Ҏ��6@�XwI�߯HY���k�Ï����j�2�cզqN\�ɉr�.���pT��~4L����WLp���������+���6��K<���\�O%%pP#�EO-`~q��e�5`�`l�짪�u�I�E��?��[Lq��F��x6� Ÿ�p��摷�2�3�	h#>bb��𭦀��?h�k�WL/�Yt�T�E���]>(�q�`�/�����=u)��Qۯn���g��6T2�5�b	]H���Fp�L�ˎ��ȱϰ�8X�Ks!Ao5�$^[�ƓQ�?��-�/�uNWϿ��T$n�����#�����뤉K���l�{�U͠�r+�O+���$����D�,;��y���L��s˧�[`i��&6�L27��Y&"���~�(C�yy�=�޿O�
Sr�\6j�D��]BGIB�E����#�H��L�@v�՝v��$q+���j�G+F3�G?�5�3_u�9��(�EM>���џ)��/W�~!�%�/�2T���xB?�`�Nd���߆�J �
�x�5�- �m0t��[����32t�,�P|�)�sC�2S��
� `gPeTɐ��Q�(y��3��'o��fԋ<<<2��f?[�k.�(7��6��-��%��t�����Ӷ���������߿�J�Ck��~�5X;O�8�����e-&{��}&'�A�)�(�����v���ڷuc�#L��Ŝ��������
�?�/�&�3pJ�N._I|9zԃ��}��`��^'�J�luwu�<!����X&g°=�w�m�:��f2�X���@�+�E�̲k�翹�hO�W3��y?R�˓����w��b���d[p=#$����l�oP��UyI	��6���0�Mʳ�߶h���D%vG]����U�$}�vPD��Q��2��e�K)�p��̆�����uL�62������''�.Ve@��s�L��࠽�Zj�f�zbb���]��_oeVb�8��mK�h��H����XA*��b���7�e�z'߁�2�����u�k};$b��[	��7x-���ybW���g���u�X�ɛ%֪��o�x�߲}{@y��4�N��?�J>ȸ�Q&;��ûa��v^�j�m�)4�/Ǎܠ�Ü�f�bcKò�|Q�!��H���nnV���C�(R����T�PfV��7Ք��4ESU�:L��"jU~���	B���{i�%Be�)��J.�ZY���=ܺř����kaG��P��3�	�V_@C?�6m��g|���w=p�ܱ����ʓ.��`���� >C�S���?6��,���,��^�� ��pZ	���b�J P���Wȅ>e�8��)��e�	��JH\��9��H=G(����b�/6��D����m���}3Z,7�
(NWR� �����r*��i��>%��~/�pG3hx�.T��ڿ+�~�;w�}����<I����Qg�x���v�As���s6ъ@h{û���"2ʥZ��MC�������3���G���ɀ��-UM���Ǜ6�j�ֈ�Q�Ci�E�Imq�l�XE%` ��]�wM�J$�>��?�E�~L[���`̋�������֋��YH+�4 ҁ���5���������(\��P�r6��� �r���5(W���۔��O� ��7@p��|�Vi-�QQ]�1�q3�;P�&�������SND���D�2v0h�:(������hR�<y�cu��p�t&���ͤ:�ڕ�&�ܧ���]b�䮁��i�]\����G_Q�h���S�o����>EI�Y �y�f��ٕ�Z�c4�������9P��b�;,��'π"�
_H#O��͚��T�e��0�:Փ��r�b��n������J��ϩ7Ct�ز�E˨0*FnsZ���r����fSTn�j6�����J������8�u��xg^
Ӊ�Y��1?�tl�@#..'�k�f����U����c���*���)z~]�������a���,��=�B���ݫdԋk.�k�����@'��`�C�?�m�U�Z���аT&E�W�ۯ�-�\Y�����2�+�J1~��V����-�gk�R��yyy�H��hQ��p  ���\�Ía�.�Iep���,���,lQ����S��e��Co(����&-�`n0��}��R�Q�X�6L��`�o��\A�Uf�Y݃e�_v�o/@�4��ɷ��~�4�7!�<	�A3��X:1gۣ�k�
�]�$R��������	~1����%�] ����%W|�����ٶo4PIq�m�%�E�����9�(�m��f �,�� �pw��+����9c�b��89q*�9��rS�2A��p�jފ����d7�Y�ދ��U�?��T|�>��~}�F��c<��Q���L���V���9߹j�%<�c�_�{v����&�t+z��Y�֯���o����΋�':&�[����'ԩ�~�T&����n)�,a�8����?���!��`��ۋ����R0fȮ��
wp��ܽN���[��J��m��ơS84V�t������3���-��3Y��A� N�K�k;h�~���<E�j���lǉ����u۝*P���=�>#�fZ�~Q&w>2�0oֵ�ã#^) !H�r���%[��c�N��|��o�I���� _C����*Sl��)nAW�߂n��?"o��J&�"��w�P�2|_�Ď��t/�E�/jR��%$S]]R\|k�� ���g���?� &^����߄{�z�5^}�����u\�d�.�{,�rMj�Sl�}��c�����Np����'��IZ`�Å�%��1�|�Bh�T����b}0'y�$�v���h�ys}1��Ǐu�o�����a���N%���d_�R��ԁ���|�$#�FgR��C1w�;�{oS�̋"���p�b[�0�U@;�E2�|��?b\�.��@�[E�i<�?wj*RAc���?�ӱ
6
���;&�@��
V"V��>�I��j�F�;��8�$�o��w���3&��)���d�]���W/�e����H$n�i�+@�~v;U�E����QbL}��x�e����������nǓ���Y)�#uC�.m����X��,�
u�!��k&1 ����#��,�9��[�<<�/x7�O/"//�ah��(�M߿=���Zn,t�Q�������CBN��UB?eI=�/LN�ozj�b�t�h}a��J��s��G�8e��w�4hQRD��hP�T�2p$u��������jKՀ��fͶ.L�>�s��m/�f�Q�c�?���Waø��?�����X\	��.���R��������F�i-N����xȘM�1.���Xc�-�X�C;�"dpأ'�ò���|Z�P����ǯ\`p�FY�I:4L��\Ͼ2��{ڵ�&Ԟ�n�VWL��^Wi���U�����͐r��E+����%�R���u�v��B�g���fsÄ��F�&�`}��R��@�Hō��3E|v�>Sr�=����#܎����4@��[s��Tɍ?�B���p�c��v���:n���>�C���fT�mH�p�b»�^]	0�񀐊W���6�x�Tq��r0�U�����G��Ey��vaU}J��j�kL����Q����/hk$��� R���߳�뙴(�Z$#��;f� 2�N���f�E	�1���O.���,C'�j�}��&n�V���ۨ���i��ߟ_�SJ:9O@ �$޹�E�|�ŀ�n�x" br �sV��\��$�?e���n��8�pDT{���*{=x��(nn	Ȣ��mZ��]�o�x���FV�t�v���|E5����W����! �0M�^0��w�ct+� �O��$�E���/���[�$��}9�������Oc4�l`�ŀyv �5�RP��[�g�8�`��ǚ�2�ֺ��g��h�wt�E'~�[=ʃ�~6$���$�����G���A5�=�Ž�[G~[���2S�D�Ȏ8i ���N���3e�K!��$D6��A�	�l� W�&��������Y�c2�	O�e��kU������|{v��:I�!$Cf�5s��*�N�z"J��Ĳ�Ѽ9�<�@�ҷ����Ɣy�� }V��`0�6���Cd���&�"Rh�08�'տ�  b����@21N�F8�45L#��:�Nf�S���=���_�x��?wiA.���[ (����]e�_ε�d�md�u��g>9��{NM�������u�6��E��->�:u� J��1f��H�������_R�d���d&��.�g�+!+3n��Dv�^���uq��y]#��J��������G�۽�}y�s^��8����|��ni�����M�_	��~o�y0�!v�:���]��0�tH����k���˟6�� ��M2P>;gT��<��C4�Q�A��P�� @��1X����Ew �1nD�W 6й����3�)���������+Louq����@���Ϳ�����+��0n;nuE�A�<��_���MoJ0C ^�Z����Jbz���Պ���Ɗ�W��ή�!.4t��ÛS�X�]��`	��o�ǔ���;]:,U�V�{�J+
L�+*���tݩ+x�+���_wQ�.�:dO�R�]��8�<*Q���-ܼ'���}ì�3�gb���*?VRz��|�_Ww�:汝4\�`��#�JH_����{9���m"N,���z`cp�*��,�=A����e�sG�f�}+b��;�|���1�5�o%%J��AU�L���	�R�Q�x�u;�W���� ��ț�BjU��0CK��!����P�J��g�k�}�SCo���:M3�=�.y2��_�6�>��#�ȟ]�s�d�ߛ�\��@I��g��C��]�pSk����Ů�������pw��[d�~�PA�C�� �e��ת��_�	,)��~�G�]t���������5٫������~�Xφ�d��f�
�@	�"�O`����?������n�ǧ{R�ߦXY���SY�����~������՜�_?���p���i׳�>�������#Ns�7��U���&��� ��7�����]�|*P;��,��"�]�w���y	��J��*^>���R�X����".8_7f䫒ϋ������
����-�qL�W���|��P�|P)�b�W�L����,G�d���zb�P��ږ��$NsI6���)��tKh��3�V�=�����F^�_cXj'f�ʒ�&?��h�mk�@w���,���{/_��!
�7�l9��2�7 P�gf�y&��A}�؝}7(�[�$@������A����a��B��5}�|3C�tJ"��ɋ����3��]���orV����Uٔm��A�Kx�&�x�'E���~M"�����#f�f]R;D?i��U���xhg޸q�$B���s��s�#.ѼA��t����dxh�n�}d5��{Ƈa.�}C�]�7�l�T��<�	XT��
t�8?{�o���";UaUqz���ML�?�W��R�3�"
�n�7)r�ӏIp�'k�S]����!�4�=L��q4�� ���y�y�����}���gj�֍������!gd ��
��?�T2���7w�����Pέ�QKgFs�ԇ/��݇�n�"x�v�w��G�m�������cA:�Y�Ԏ�(��Y�N���gײ���Q# *	��(�%����C�M#F��m ����?i�vaE��Mvˇ��j5�����H���7thŠƵŞ��T���T�C��� �7nRq��$|�n�'Q����*�ض�(|��]��q�J�1m�S�*�d^�� $m�ͩ��,�e?¿{�:�2l���#O�&@��ʤ�Z@�$\���nDEѧ��0keV-{�%۬û�o���|�Q��U:2�B?�v��yS���b�=D���~�Psq�P0	�}y]Q��"�fP�A��a����%n���t��L�
�lj&�̹�

�u�3σA�6��o9�40���Z�lߙ>,���{x���a�L��TRu��F�m$��c2��ECC �0�9 ���i;�����ͽ���\ߏS�'����9�E�`�dr:���(���oЊ��Y��{n��)<%���	�{{z�} @���T��'��?XUY|�Y�Ǜ3�>��~�l���K��(f�����H�i
�]��+_�E�v�m_����T p������Zz��*D�R�vviV��q�.M�n������W��9��õ �"7�ce�k���rǾ�)u��|3A�tf���r8��J�F��L�e�!�6�{W���؎�ǂ�{��bUr��4�9 �1�xh!����G��lB�ٗ�PV�..��r!���n�*��X�+���
?�Jp�d�� N������f�/,K���.��f�����\\S���7����T�����s^ݣ�=�ZDZZav�m�,��Y~��S-{�/�a�f-Cf�-�W롶��na��o�����B�:Q���N#Y @Ƕ];��gY�H$���AڬW���!a��Q��e.�B|pȗ���y���<���K���3E�;-��N�i=��E#0^ёX�l>�7+��ao�9ģn(��pS���U�8R��)�Z�����?%В>qy���]Q�:�X-�Y���з�c����z�����G���{h���u�ę�G��tx	}��|��(�/�?�}wZ\���m�
ƑQL#�R�l{���=$�O�qK��О��;9o�y��Qn���Q^�t��DH�3����J�0�m�ۂm�1�|����_��5�R�PG����"���=�=�������Ұ�|�a[@35��#�A�����ުO�C�Ðp���z��\Rh��mz˦�dϾ�(rcF��s{�h�#7��\��Q����y~�7+�.k9����P1ʟ���o�j�׫)9�WJ�X���?�?�S�]�7���/f�|���w.�'O��u�p_QT���&�L�����c�y�:���Xy�F�M,������荇3�D��W��I>����iv>=��_/H+��yc�}��Է]|�p�����/&�|�ԙn{g�ʐ*�J�<�8F����n�HE�q�JH����Šg�Amb'X�'!S�	-�������?M8TY�y��=4do���/���^Z�og�#Pu�O����E�zYmj��ʓqE�	5D�"'�A�H�Ot�8����(K�*2�8��|=�-i}q~fp� �`Ԫ�9�eyS�b���{
FCb�Ѧ��	��=V�\���k�N�˓��Q_�
�&a�Gꢷ;�������:)�����ﰒ�.������|��n���)���ެ�q/!��3Q~���/��W���$?�ȠJ�hh@��$vRl���t���}�J%�:E��t��B�|1&�a�'k�R"8n9!�W��R=�*���S�ua�>�+!�&���^]Ơ�9��8�7z���[9f�[_5t[�;|EZ���ҷ�5K6��]�/�4�@b���(�y]F�`Րc�9�@�Q�n]��c�8qԣѭ.óR��a�q�ߚJ�L���م��~w��J=9�GV��c�4Ls�	��h��xƏ���OPOަ�8�p�7�K�3��<�}:�p�Z8s�!�V��q;�H�
ަ��<c6����[~���� ���V��c���#)fTn�x_î����t'N���}9<������P�d�z7�e
��k��n����ޫ2P��X^%���*��7i��+�Q�T᧐#Eլ`y����P*[�� ΑG���⟽́qZcɡof�7�SM5����c��o��ǘz�s`0�Y�>f�:�����m"#\�=L+�&��l��5�Vj����ʚ������}cU�oό�a�υ*J<a(��5MXy;��h������~��4êS�عwsʚۯ���&�G�����|t%���.9�F��44O�00�N��R��H��Kq&�ɗ)�q��a29�I5� Î5�IM�)���H�bS ��*qX~��C�6xM�/p��j�V'p�����-�;-1�"y�dS~�Z%���$rv�[�I�@�*%	Q���	2���ě���~ic�f�C>R��>�կ���LsP�P���}��n�BqW+��d_Q'a}�TN�n��ƨ/$C��C�b�xФ�j>�=�_DB�#`~j&�Ψ��F�g�X�_�7a	�]�v�/���{ݡ|����Z��*6 �H(6 ��������-LrrrC�4�4��a����Xޓ:�	�4�n��{t�axK�ڕ�c/u��DF;è������o���$DaJ�d|��_������ː�L����-��c�R�V��b���&&!g"�1����ߠ7�.e�����Y :�!�:�M�(�[I/t��y L�>�����[`19�y� �/q���q�(9�; ~�۴o0���r 3oq(�qk��gSVK�_v�}a~�����J}t����j`}	g̞I�y�8���P���J[�{t�H��'���9Q�!���E�Pk�����v�F��鏆��V5]	�G����pK�xʄ^��Q9!����C���?��_��;)���xB�#UT�ˤ�p�%���7Or�N�;pb00�G�y.H�_E�s�Pp%���a��u�G�� �:�j=�z�����^VV�n����1V5��׆��f���Z��*O�_�X�w;�J�g��Ci����}O��FG�CtMG��bS�.*A6�e���/��Q�����V*��J�eT���b��[Ӯ�߃� �5c�}u}iIx��=�z����3>ڭ���j/�wC4=\$��w�do�o"hf�6�a}'����c�m ��t��������R�^´7
�?��T�<��[��\�XiH�22�K���2�D�o-��ts�Uݜd}2!V��(.F$`m*I��H�MQ��!!
�g���S�TB�f�%�A���v\��c��6�ҕ��^#|lH�>.ɘ�&J���:�07��Yr���i�>�$������ (����e�
{;dFW�T��j�qqv8��Y����:�5�|؛��7����5�gC���sƈ�^֊����ݣ�z�k�6�_~�����UK�,.%�w�� ���U�8:�S�z�w��!�L:EF��#���#�0�]%�!��2���ܬVF:gDde�}+�5�督�	 r���1o��z���q ��?��ٽ�YQÙ�hO��j�m���O���NVA�dDa�C��Ɩ�D}DkY������=n[.G��r�It�Ԡܖ~�̣�k�U�q&~V�+ؓ^�5A�� X ��lv�o�~H;x�6+�|}SE�$��3�S�b���F̺�"�d�dBy��K8�g�fr2y��[wqn���|��m�V���&�2�"�������[�06�'��W�k@�FҘS:/�e�H��f99k窿���ƣ�������TXܼ�>jJ[`���T��|�/����m �<�M*D�Ƽ�rv�J��/�����,�v$�f���N�z%Nr*h�))��^9�$�(9�c�P�p�:��ש���㞫_F�5�<�;%g��e�{mHi��MT�S���		��/.V|J��z�މ1fSp��cg���������0�A�;��<�M����;��I���l�4��iV�3 v��J�{a�e¥oN�I}3kh��Cť�l���^e�=�y�vk��9]Q��.D��a��L�����v¹�u(�+e2�U���&��<4�N�%��o�Ѭpg[���L��fu<N�,�4�w0%��a��"�W3%�{���w�}Cq����vA<	ӑ<��z3-׆U���R��Zr�S$��^��o3Udx�xݞ�����>�d������rB}S
�me��L��8F�
��f�ٖ ����ᝇ�"J��@��#�դ�u���?����n}���T7��;X���Xl8O�?Jp3�k���儚�"�<�3А�����y�Gn�Ӄ�N𸖶���Xu���iC��oEؘ�ϥ���-T�H���V�~�!&�^��yW��J�z,��IY��B��-��K��S#c�xL/�aKN��s��7�@�'��9��f���a��`�XR�J���<�/.?��"��Ar�eS�?[z	�99���p�{ф�#Ħ�`��>3Ʃ��oR�jy��D�ơ�K $2B������3���5���}!�{����t8������)��!ύ��?�3��P�� Л�r-/��z������ wV��Δ$s������y&wqP�Z5�ye���/�:8��˟Ύ��iqww�LO�ц}���	'b�$�	��ɴ�1����y����÷_H
@��?��[jz_�3ұ{�X)�-%A�� '�$��5��0��I�����5�::p&Ü޿��C'�U�i�NV������% 9b��,D��u��~+�ֻGd9�[buvC����i�Q�oޛ��q �f
t�0`��k���I�q)� ��t\��ޗ�r/2m��7J^�z1��[�:�w(k �gݙ��o�R��"L蝏5������pP�� �$О��!MOJF0�H��˂��I0r�y���*��_R%���?��L�}���L�pB�ř����I�)l	\����6w��!�t-N��.Ɣ[��	g�2l;	o�r�Qe�%ab�[bO~p��B�<;uѳ"���2��xq��بl��,���7�+����~���K�(_��x
/����!mV���%�(2�>�eXG���fT�lP�_�%�nꁻ��Y�Z�P��?r�s��]5ǈ)���i��{WFLEB$�D����Y����:3Xh���R�Y�I��.�JYF>-���[��m����qP�~�oNI@x�7�zN7�*ԩy��V>��z���Ez�A%MSBo��#�w��#X���*A���m��.���a�׆�����4�"�,S;���ջ3��������d=Ȱ
���h�X�ٛњD&u��'�h	=6N��k�K���:���4�&���1N�V����H�RL�>
��z{+�����_�(o�i�c->�1��F�y����o�(��@���8u���-��=���ϛ�-�x����v��F�q����p�L�t���Ec��<���zz��i�I06�#��a���m��	p�9r����fS�ukR }��T�e��J��<L��V_z!ˇ_�dfZқ�Y� �#�un�ॎR��o�o6�_.o�Sa�ɫmuR�L|�o?�98�'M�z����<�������|��FՌ��҅1/�:�H�й���O"�/g��c���+�Q4������ �a��&�+Z1��ز�2�~��c�ƀ�����5)�C�ՠe�����莈��㚅P:	��;N��Ds(��Q�\e���;���_�d�u*��JW?��c�G;�/w8�4X�/��U�ov�Q��r�� �������D�;_�f�w�_<t r}����{j���V�z��t�$�#|���,V3b��sxw^���ڟ:�4U~U���'�����?�u�K�Q_[��<"�?�"^�?�����u5����/��d�����r�H�vj��?g�\ǩ��˭�YѡԘ�nu�;��H�J�v:���K�?�j�ٗ��*w`�=�ӹC�����wQ�#�<��ti[�xx����%CL�����h4R>�̼.c�������+'���_:���O� �y���5�>å��1����C�Dsk����-�KM�WC"��|�v5;�M�e�Q�� �(]�E�����#�^���,44�j>s�йKG��Ƶ�.����VJ=��a:�z�iE�1O�6yPI� Xw�R��a���m�KW2�a'�J�i)cu�e����J��J�E{P/�R�Vg�}8}Í)vsgBZ˞�r(�sX,H�I;�7^oO�^��V�����7$D�=T�Jd�rk�"��g��ω��$��๯������B���n��q�%�Hm��ᤧ9]������h����y�������Nt1S�2)���%D�;T�%T����~u�F��i�}�
��v]�v:�G���K���I��]T4&���{_���	��2`����qD_��6�9"U��[���i�����2M��ۂL�M&���@�V��N����@��}�a�\��/�r�C�����6�g�Q�s]�{d�,�I���x-(��L�!4�ZoD��<Jdyι��햒R�A�m�3aIބ���U���|��>)���xc))�s���QY���U�:����z�G�ĵ���<�3k�J�1�Pql#�-){)t�:/���f�({e`$��6|@�fH�j������S|��`;}��f�S�`��"��i�}+_tsIÎ	 ����j'�g�3�H5��IۧHroO$]��[b�_N�g5<}�3cT�J�����w��?�n?گ�K�������96?Q"\E��(j��Å%��Ẍ́C!	xbb]Pq8���������+W������'�T�=�)�bU�Q�B4)�oA�v�h�����ib�$����oE��ŋǒڹ���;qMr�������=�_'~��8��w��m�
N�(����H����lҷ15�MNo�ȭ,ed�R�P�&T�ӝVv���4
�g�n �&���1�S�����R�Y��DV
>7F/ѫ���Ar`���(#�Zl���z���@Ô������a�q80M*�>�����0XB�vGj�C�3����nvC��N����'��'�g�'��)I�&��.�gJ��M�;��}|�[�uD�����,�=��&^�FܘbN����#2���m��B6�)����3���sd;�R�[������G��*K�g97�O�6�f�����#�yf80�O^�8��v@�!0���,���6�L��- >M��Gp�0"�MG?c�{�TxHE�I� I#e��^�����MvX��:h�KBFT6��d��vɘY�?��Pr!��+K��~�_nO蟭��E�����_&�Y؛p�I����?��t�=�)X�.N�.������wS+eyC�B���� ��	S��Y�N���6����Ҝ��KO����T �qǡ��?�����a"�0�
���_h�|5�/�7�H�q��Gkx�a5�C�����}�1�0Sj'" ����G�2�$�vx�\�R&�%E�L!׊u���I���w��Ͷ/�&���s�jjY�����/�5�"`��woXR�9+2v���C��<U$��t	�+/�咰5)�Y� F��&����x>�� XNm��4!䐚)�yz������D��:�mɻC�@��!�Y��t@�m���#1.�G�-�X%%��>U�����Q�>m�����ie��}�ר���+��G�+ҞV�}egON�����2Hr���Ws�����K�v;���y��0���} o�.m��,�9���b�FFZ뿵�G�
ѷ��ƽ����!��r-����Ԓ��GT�lk�U8g�h���U�z��iIoQZq%ڥ���&4Mu�]�Y�j,35�Dp��|^�J�ܤMu�}��K�y���a���2I{�1�%�,�s��nN����%M��$ǧ3]�[%�x%*?�:�*��X�LÖP.�>���X��oD���9���.�ًj������2'L���V�t�Q��-�|VNH�.�l��YG�Hx��3���b��a�9��߃����o�؀�OMp��-#H�d����}f�?_� q�M �mlo�*���J��(����>+��䥫��z�ݼ9i����_AAA�����H�ʇ�+���W=�P���(���G=^�&/�*A3OV\BkF�d�+�F>�V`�M:���W &���`!��^���Ҙ��(��?���H��?�%�i��[��O��������#�y�\�&�X�	|w�|x7�M�"p�D��=Ԋ-#������l��Ցc����!�K<�Pt!$�x��~�ng���9�ź���v�ra?��}�]��=Zzw4� ok�A餌(A�e-7߰�ڽ�`�C���b]"�#`^,׉�#/]��j&�9%B,.�@��^�4}�25����o�r�����I3���c~xM����Fm����߉kw*ݒw.o�Ad�!<��,N���~��-gw��]Ȫ����#_����ƻ��$T�~��[8�3�+:��Y����T���j����[o�E�7����v�@��t��o
��ǨS���k5��%3�%Jz�鏋+�r�dڅ�*����z���r $Μ�0}L�G�d�b����(�
 k؁J�&�~5r ��Ngu�qc�X���N��^��Y���]�G�{hEw�s����ޝ��h�i+���5 j��(�x;�bQ� z#/2�\4��pp��Z�3K
yNX]���+��������ᕞ�Tgw'��D%'�T;�O�)��j�0[��Cn�O�K'o��h�M�����P�+$����`�*�����.P�.�9�~dLػKO/%�њ<�<Dl"I69�kS8b�`%�F~�o�#�y"�O�0��g��!� 㗞Y9�vlu��SR�����}k��>�=\Y�ᠬ��K<J�:!o��_�t���L�o���`�u�7�|C'�2���L��
a�*�����)x*U����M��>�0g@M&�7SIUk�T�������!%_�V�Q.��A��h�hO�NL������v��M���Ӿ�����v�﯊=�4�b�7g�M"׊�խ�P���`�����LUu���N�������2��r!�ˇ��?-`��<��C��o���������h��7�;)�Й�ZZ�-w��V�/��.���<���i��,54s��؀Aҵ4�]� t����� ���n�S$B�sR�F�^�������8|�/�3<୘�y����}�?Ad����#�>�ս%ܰJ��4;�{߶%��eO���u���L��I3>XC���`�ܮ�lҁ9��H�^?Ք��;�x�'֑[��O�����!K{����}�uH�Lw���n��42�wi�o&���a��ܜ�sj���m����nrN��=��HYlmd[ˊ3�v��Df-7��ۆ*G��w[;l��A=U��+��Z�L7Ef]L��
�ǐDv��]-=�tt�{���w������ބ��t%�h�gH��34�������	>l\4��nc��!1)EU��0g�ܴ����b�7'%����ܟz�B�δ�d1���*-��7:/�'�N��Go�3<�'��^
��a]d'����r����Yj���ר�$�`"C$���
X�g��[wҗ.����$�yN�v.��nuK{�ո)�T��(t� �~���(�* �`�Ą�`�TU�m [����L
�|����D����T�m��[��,���m�A&�Տ�Z�и�������x#�շ�+� ��#�uFJ�v?�
D���N��:�`H*{d��ٽ��-y�Z���ϖĿ�1�<�������-�WW\��$D�(���u��H��_oΊQ��z���?otڙ+\^�L_)�������1y�SVv1��
>�x�jJh}�o�K!cy
�G?�t�G+?�L�F��N>����X�З��~~�ܱ{?w���$  u�����p�Ν�Ε�;�$zQd�"z��T$D��6)^O$�C�iJ��~�'z���W)�P��RETځ ��7�ر,B��.?�������B�1ݜ��C��|��t]�����W(�����F������"�u��h���f�t
���#~^$o�������b$W44,V����hz?z<��H�;�}eو�=���^�%��8�0��F�J2�<i@�w~��J��eF��l�}Vp��g�z4��h$���E�\��uX�i��.K�![�����9v�hf҆��P�>���������+.�_����Eoa�8Օ'����Z3�L��*/G`^�������`��*�ߪ�~�,��Ŏhj����_��;n�B�FJ�;����3e�3=��k�,��"�%�py�s\6ԭD1�~�S;���,���:M��oz):��(B��p�1�p}]��_�wC�>'��n�1�K�>��Z�Z�@����1�ɞ�gKl}���3~��2�dv2L�]1�W�4/���|�G9큸���M�3:�&.,�#���f�iNJ1�,����x��7���l+�;ʄ�V���n����iδ�t�35u�%��T�d'Z�&�%iʓ=�JH�"ʒ�K+���@B}lQm9���!M����e�>⋋���2Y��5��'����-���y6K�@���&���	~��0[g�^mIp_�,��o�Σ����}�2v��F\�QLR�I��.�jWR���������@��p�r+p�Nz�g�Wߪ�{�� �ѻH�U��\3�P?�y�e��햱��a9�:�g�|�jO�oGp� $9d����>�aq5i|�7~PK��~� b�'�~��73�I`��ު�Q393^3�ݺhU'��Ҩ���0p)�%�z�؏��m?7 �P������t��B|�N����>fxr?�:'����^ͭ�Cr�KE-�-�s�t� �>߂�E��KQ��機c�y��2���P���(�Iܓp�OZqJn���A��!���[���A��E�/e�|��U4U�V�ۍ�����)P]�!�6
��0z��=_�ߴ�� �͂CZ��\2��Q��?�� �Ϲ��,�7��P�%ة�>�'���i��Ьf,օ���J�5	�RO�`������i��
�
�@іE2I�ޑ�4�,(�"�l�704�?9�X�^t���T�?��s��m)�Pa�Wֻc&�Y˯Q�kVf�^���ȥD���R�fu><��"[�V�?�(ߟ�K5���A<H����fg�f^�i_:���-x�iBk7�=R/�����%3_���пo_ن~�ٰ�����+�vq_J��o?J���Q�q��Ww|˧	;1����/�(iH�<p�Vg�F����f��������$�X_1n=�;?ξ`*.��_ �&�KE���"D�M��mŵ����&z�� @f>0���^���ITK����'jr����!�QΡS��N'�z6�4Eϐ�-�w|�!�`���3���ځ6`��6��N�h�d�W���^;�`
�{L@"�����a�K��w���=�v����>�v������d���q�k����и��,1!٧H;���n}�쳁�7��H�^�3ӲVY/W��!స;���o��j�F�ȯ���CVU���1y������%1k��,�����0�xz����	1 ӐN�Ij�I<����9^�R��/�D�cId=|eX��ڴʤj�Y���W`��܅ű~X��"�S�}� &�k���U��
<�M��{!�Ѥ�r��x�6����}[������ xfӷ�Rʇ�ҕ��r�����r�2N�Ob�X�]y:ѿ�c�g�l�y�����������
/2SR�hE�p�d���᷎��0㝇�U	������~������	��T�cߍ�H
`�6:<��yL���CIs�|)���q�����{�����
YO�t�c�(����f���� � �`�����oS������UdH���I�h<�+ӗ2��t|�l��!���#=ׂ���K+bX|��@;V�&}R��9R�ݬ��'>������5`&#rmk0>�o�Ʋ��s��"��,|��'�7T�X�[�	�ZC#��sm��z")B��,<�$���=B�Di�|b��8C2�`��W���c�U�i)�j�A�����JaJ	Ee&�}�'"�	F�+�����&��
>�Kj:	�����*A��w��& ɤ�;o���1ᕻ�r'3e�c4�g�^��0|����i⮅װx g{�ĮC���L{�x�o�6��l,��R�\�� ��Oc+��n��K�#�06���"kT��ƃ��v���]JUѐ�����@�������˽��9X��C;���~��騖��dߺ�0<4��`���f��T��KΤ�����	�Cȥ ����<fK���:�kθ_�2�(��rS�t m`ˣ�?2!8�7p��x�`�P����a�V�������H#W>�9^�<��0cv�B�8�Z�z/�6ݢ�&cD�Pc��e�v��A�<�����)�������3���ozC�)t�x�),ǁ�0����j�9����ي2����2��57+�/6����XN7zVd�'�X�J��Vvd�W�w�)�z���o���p�X�\���(F������:�A�����;��j>���=��]&u�����q;dU���j t���G����*m�o��0��d�播�P��B>�8X���0;:Ӓ�E�mN�1���h�������������3>�4k!�NV�����<b��vs|}7I<�e~��_W�𦴇mn���(����a��X]s�Q�np����=6�M_�@���?`���`w��)�W��	�bbrl	hN,IY�W�����Z�j/�����#��ŎCa�&Bn��0����@d�:66�]���V�C������kNnn'�%X�� ��k�U_����t�vu]�)%E�+P �G�_�ގU�8��U\�$ �n�Vm��=ԓ�w���ꬠ�fU=WA�FU�@�,����0��w�B�{����S������ˬ�6����ZQ�t���N�ǋ=�v9R�/+B�՗��p���!�W��5��T�	}X�pu�˻w���4gS�����(B^:��	?2�i9=��xK���7�Tss�v2���]��½0/+�lW��󕆊��2�u�,'�/�����_���3�ʏ����Q�č}���?-�[��3�rrr�B�.ӾSb�G0� }��[G�^v!�&�6�޾a�bs���w�� �3W�!٠������Vi�C�������ܚ}R���_����rN� U>�V�"7:�Om֒ON���I_�:\8�����9��?�������)kx�1����O�,��{{k��+c��^-N�V5�����oN�j���������|W�t/m�佢�ϯ���)��ɦA������T �ɚz��}�.ښ��0�Ή��}�
@��7�*A���Ak��K��S0��aBR{,#�_k�PM�Ջ;>�(dy������ϳ'��^�|�<��&��������,����p�5��C�srMank�j���A�����mB�;�&�h?�����ѿ��C���
��)o�������펑oh~�2H+];eS������� ���&�!��լ.�J�w�� �?t��f%�Ѣ�)Y�9w�w�7�u���ks� O�<,<��v��I�����w�m����!��p���Xכ�S5'�o5��PKUw��u��\;�&O��/�t׉�PoـJ�6�~�+��aနTBy�b[Z�� _�׆�U>`�|d<Q/E���xL�ԸS�(�)紐�1Ы ؔ��]�;&��!��L���&a��JțNh���b�˥������C�Eڠ��"ۚN����(2f�&)0,�P���B��W=߷~&��u��/VI��e���B�tC�R$F�u�����{2�M)��uG����q>@&�j=v��v?$�_�9���G�Ҍ�O�q�"9ti�'UO@��{��{"�d�>�����2ux4=hj8�|M��ù�1$ϾO��6��X+�@gF�3
r
_�t��{~�vtqѪ�E���%������c���d=�2r��Q�u����Q1g�J�j!��O���JV�dt�Zb9I7x�M��Y��s�����:�6)j����3eu�G�i�W|��C�AE> �����	�.G�CGN�W�4e/3�e�m9u0�<�)������C����}uPo�y�!�X�L20�EN~� ��� =k&�M�!��b)�ɂ�#h`�����o����V,K�'(�?tk�7څד�L�ȱ�����t��/��o��Ȼ���G�9��`C/~kl�$a`.椇��Ծ�-t��z��lò����U�7�⹌�PKġ���ύ�ʘ���c,�~2��*�9m-�.V�A\It,~�'������29!h28x_�*˃��}V�V�1Hv�ϤDJ�S��Y�)��_�R�P��8T��8�$����ce��.F\��=x�9�Or6�n��{3k�?�Z�e�_]�!�������L�8��=0Gv\k�Y��N��{�"��N|J��=dl���F}���g4�����7�3#"l<-�R���7���NF,jY|��?�ײ'�B��,ɂ'��/G,�����~�w%����!���_��J F)(%Y���nV���YIGl�U���%gi�m#W�`�nHܶs��]Qsl
���;���_ѕ�q��"c�+�;H�sb�|��{����Sp�q Z�z.}������&o�T�T6(�ʩ>%i:<�p̨�D��>���y츞��ݰxXe�OY��xbu����i��e$Ϳ�����)��~�H���C���pW�����Q��l�q�+���o�W8�dz�=�T�:>�x����~�����
���#/�K�rS$�����.����G=!,.��Ǚ�1�6?�B�,I٦��Z2���"��&�rs�f<�W�kqaI����t�L{� *"������3����3��e�އW���^�L��t�#;��*-8��s�D�A��M])ʝ�+?���`�^�O�~��W��x�6�r{���!G�ڼ��MU��.�!�|�}��?8�mF�ާ�'��W�QO�^�t�X��B�댆��plv�w)��`�u"%ս�g��U%>R�
Ǣ��U׹P��_�.�#�g�U�%i�����:7˄X�]|����[�~FoS�R�6r��z2:6�B��S�%*8��ĝ7�(]놗���N?<Q�=�N'�tz� R�}�bѾ���,���h�ڗ�"�@X1�B頽�dE�A�P9z}�m�+�`�i��Iܳ��~�Z(t��N0\��g^�ߞș�vq'Rp�:ď��"fO��'v��N����hoD�b�C�r�H���HG|y��_���-���e�����.�FN{�.�S_�E�>�z��5ݶ��w���%��O���恤�A���d��̆cH|�t�^k��J�+`S=�2�pV~vN���+��4K�V�d�+�[Lj�cUO���ϸ�{�����k)��K_��Ɓ�2H����[�D��S)�+�¶`w&��]��������� k�{�@PA�7�*M����Bo"% UzQA��� *M�tH�"5�H�H���N����w���!�&Y��sf����{2����Ss�3��n��X���{tT���}�5�eV�}
����k<���ρ�B�s����<r}�O�{�*E��;�f'y7�*��o�/w�!lI��h⭱"��������J���Ҍ�g�Woj5�[J�=mv?����1b��E�J�����]7��Oi�����DH=#X����Aڈ2���K�&F��w�h
�3��l^J唬N����U,�=��#AfZ�Y̾�+?9����i��r��M:E?Al}�PgI� >U���9߲��B�I!��~� ����y���+������^�a��C�J���B^UTT�"��BR /�Y���p
�JWt�4"�ocSz���b��_����(o�>��ԋ)/�Y�7���ۂ�] $C�0�p.���:�}\�:sZ�n��\�^�rn �g}Q�'A���;�ƴ8{�^MP�$��%h�V&b&q�̛}T8TCC]]r0����㶴�
����%�&?�x��a�K����Y���������d��Q^a_�	�2�M8�-���i���;wZmj�&!B �M��cɷ���\3�_���0D�X:���\`蕗�ϬI�\	���i"g�T~���C�Rz�v_�'��
0}re���$���p�ؠ��Ѣ�&�Ĥ��H1|�9_��� \P�*"G�^�6�X����EԺ����߸r����4hx��5)]RE�<��*{�x߳��fE�8���Cl�W=ҳ�c�y�/�s<��h���=��k4%��kYj��m�m��#�r����E7���v<�6j�J)��I 
˨s�9>�t�L����
�u��锚�x� F��M�P�� ���H�v/�b�� TV�bhѱ�Ҹ��"�v4�[=O�Y��2u_:+P�?��5u�o��x�Ue���&jS��B�Yi�b�Ͽ�����&�LE:������+��j����O�Ը;rǐ�~,n���Q%|�59�愺�Pإk}LPh�u��*�xr�w>�˰�v��vq�e�@V>��y^Q�����<`Y4������N��V��)o��Oh�r����\��]����g'pP��41y�\Z�[롟� 'w8�{����,� G�-� ɌT�p~ %�߸�C��O���8�|	��}�=��?xv��#���>B��Ws��-��+�	k��Y��	��!�髩��Up�Y�o-�i���� fk/��S�β�U��������f�2Β��y@�A�d�Be�s�+��%��CР���o:��Ċ_3��{�ī_AMw�t�U��N9jV��]���،f�x��)=><x=�F�2�|Y~�S���K������bڂ���Z��fo���k�r֩`��R�N�4W{wؕ�*^?��Rқ�PdT�Z�8g϶7��LVңt)��!��
S�Ŭr�Ju9��u���?�9�d�g �\(���xW����]��\�4��C�!�w�$։Ïk�����ƕλ�9�鐬%���Ȋ���
������t�	f��D��\���ISK��.=}��R��Nk���Ǘ��y&�Fǣ�S����{�at+}�-</�&,�Z����pZy�קG�%�����4n��I����y�g��pܪ���'�E��:�9؝��D���U�������:�nsKW�V����b�q�y�_��� �(������B���qi�?8}_��4�M��"�p��0�A쨹F�1\`,��⭎�Ac��ߒ�8r	F�"OG����y��b��o'a�?X�K�ۤ���Y�A�gs�;>u�[�(z���yNj����p�(�l�͑�wD��A�?O��T��c��]�e�Q� "�� �CNr��`��r�ݽ��J�O�C�M��}T]�+x�)��{l������X�>�G�/�|��`� �9�EbX��݂�y=���#�G��K��^�	&dg�)�Yv��]��i��x�Smh�����<W�=�O��NS'97 �|d�UO��JL.ڕ�ƒ�.EE��U��xlUVQ�z�"� �g���(��-���V����|��&������X�!5�	���qvQ������b������;���c޹��g����h�|g�JF�����RL&�ۈ{c�u��uu����L��
�p�����mj��Iv1��G�ǽ0z(&���~��q�U��DKk��EJ{x���zP�]�°��v��BVv�']�pAF�U}F�*#�4*SҸ��n�Y�g��EL ������-���a��z�`����.~� ���1�d�;}':r �1EV�	�$��T]�5�(��I�Fe��a%�V��Y␼+��f� �El���t��0��q�p�x핾����-�Ƀ���B��c��'"���}!J!7��D��ݣ�a�L�vf���]V~��G<(ox��N�N|I�A�8�/�'���drJ"0!H���"bW�р�v��O[����b�d�z��M�z��U���:����0}��}r�|���؞V�x���o.�C*ѳ?0�7�=��1�x�J ���3% cgd��m0}��CO��u���>W��� N�}��R&�$�@���o.�q}O���U[������;�z�^�����z�	����`�<��⋈�H�a�_9����.�i�m�V�1XB�*
�<o!����`s�}���w�/��V��F~�����)w����1��w�(?�	^���<��ѧ�-X�gN��]�%�Ϧ0��˴�Զ ,��ˈ2�Ɂ�6�� m�漾(Ὢ˯ �8U�k7�p�ywև��K�U�my�A���Z�nw�gnnn2��m����"k$�
��e:�K�E��}R
��b�񨘛�"�)����J�I�\lܼ0O�z�����m(�\� �{�U �+�oX�����xf��e_W�/�ͳ�E}���:�M�;�Ĵ{�/�f�
��H��a6�v��T[� �;��l�զ��P� ���,2
����j�.{�0��l$d����;f�ϓ��I��ټ�W�#�W�Q�4�8�]�/Y&��r��Gs��c��S�o��㆝{ӝ�"�~�C�sKe�*�>A�$�+}�vp;D ���0(���k0�Ȩ�w-���=.\��\['��^�It�O�,��Þ}z�ߘO1�r?���,*b�W1W ��c�'��	G��)p�L����u��ofj[�i�m�/ǋ��uё�͛�R�21R#���g�cz��Yn��&�j�=�=�a�E��qx19V���,s��	>��=� ���[�kW���^�k�U2�'FѼ��n�����km�?+'��1$����GTzT5.	�9����v7� ���F��g�Y�BD��������ǷSo�*�A$銊k[2䫱��yeH]����X �7O�����˒ y�駸��\�'q����V؛$|7�l�ۖ�F�����$�-��Kz�*���"�Q)>TTT�Z��_�ng�l��Cw��=� ���ԍ]'9����|��2r�+�ɳ��!����V�*�ݷ�w>���LD�����=��n����^��Q���V�"^۾~�"�"M�K�Uh�f;���	��j�P"*�97�.s���r������p��k��L��pɰ���jה����6)��j���oYڜo���� �������i=S�g�.� ��L�i��B�3lWWY��xi\�LA�1x�������O���=�e����]<�t �Pd��s?�K��Ze2]���*O6�!��'�m\���m�?��&��}�������P*;��U�GD����}/��o�N�����=i׎��}���-�GȷSB�wGʀ`S�H���昮�l��6l3-�qe/����͑��I��z�tm�%KnP���
�sJӧ'$��}��S%i=�*Rs���Ywr !>ؔ�.R��nt\q��󎁖bi��[c�Ғ��F�\��7ߖFG�&�۶&H�����@,~�Qk��?R%;p�Z�����g������rV0Tb۔��KoU~-ה��ûHա�7�~v�Ϭ�Mvd#E��= ;�5V��Z�(���G�W�������{��{�⮿8�.���?�(�Rw�R�Z��[،��tZs͝G>�Ǘ_�n>:|����H�_t��M��B�n�eG}����1�Rąh��V�E{�~�dݢ.�wU�>�֜Q�''~���0�wۡX����`�]�=|���ܻ��y��_����D+��u?��P���\5_����$~x�kk��y��άBZ�Fe*��m�B�Mi�6�HE��[	�:O����0��N�c�}e�a4�g^lg�z�3������q���n�����&�訩O�nS5�j�f��mpE{YG���IG�vw<B�z/N�>:4�c�f>K���S�vX�sZ��HD����3S�[K�}�@,��4����9��5g���w�͡/���� .�l���p�<d�V-pFM^}�{���d����j5�Dc����е�5ٚ���wc=�����|�ߎq^�g�;����c,�I��>���R�5��CL/�'>���m������2c����̦�̲���X������nwj.F�+���k��3��FX�N�Wm�Z�_�"xlUz���*D2O���.��%64Ԭ��\[��<�"4gHV�$��w3�/����#����d�TC����~%v7ӟ���3���*�ʃ�3q.�HN^�DZUȔg.�ik\m
�LP��9yH�q��j*GJ��;��g+�|�)�G-��A�k-U�E/N,�+�oU���,���N��9e?X<�|12�Cb�t�N�e�lb8�w>�W�U��7鶾�J	A0|h��O�><���Xb�Y?�5�V�b	��wR	�g�a���*뻥�^��d��}/)1
Y�ԧ >N����|!���gBH7?<�M�ל�-��m<��M9��FJ���/iN�g4�?"Ñwp\��_�S%�>=���:�@���Jn��B`���1_n~(%<X��-���|lͨ� ��H��^�]����B:��L�I}�zvm�S��WaA����S٭�/j`�4��ǶND�.�����D��Ow��̗�i� �ă�:L*{a��>(��
Q�v*�����=���k>S�y�.���( x7V���>˼ꈊu�<�j9���)z�C(���as���ۯ�Y�$�S�*�t>��xx�f�����M���?�R���{�"I� �4ԔOY?8r�T'	��82�\���{���\���}����w�r��c�"�����q���l2!�S�t�듟���͂���7ۂO�%b��Ғ��>�ώQ]^���WXT���g��J��f:$������-M��	���R��`��[r^��t�Z*U�$U�wb�?�	K}�X%�+���u�	�2�a��Iڂ�Ϩ.�|�#�w��fْ�_l���d�����67��|��Ż��w�P!+��|�k�j�t+�y�O+�`Rj�U#���mf]�֢]�`���}A��ÐK�~�m^W��_�7~����˕�]4��$;����(C.$>�[X�A�;���S�lҞ����������c�c-f)�Rg��ot���I1��7��@2�h�>�'@����^��2��8o��sqf
��~T�.dJG���p�Alt>iDGMF�(� ����9vo�W��Hh��␶?��SIQ�d'y-LQ5oMh�"�O��=�l4X����%�V�S�[ޑ�[/�0�� ���ρ>�?G��ͫ������
߇-�)y�gx+L��=[��J��,��w�4�wS���,�|�ї⤾l��&��*���D��^�N� �^*����d����2���c{ץQ<�&��P�C�g�ت�]�s��4�`� �?噿���Ƙ�&�~u�z��d���<l��$���?��'���_)��2�C���`}xn�i�������s�.8����B�Aʊn��><u�v�����Q^!I�Q�F�Ӳ �(sH�+W���[éƚ�e�J$�"�� ���Ag3:PujC��Ѿ �)յ*���a�B���Λ7�K�ȖJ�Ϭ��X��ᚹnFl4�&D9�{���G��7פ��D�i]�+�~�W �L� 6����R �p��C��z�Qsv<=�� � B5r���4�]�*q.Nv�5J�hj���B�i�ǝ�m(%	��g��|����Y2��.#�6�){�Y@f:?t��1]��'E����I�p��ݍ>~\O?��ي`L��׫�ΊV�֨��O9��Z�]�;�t����:��J��	����x:�����a�T���[��n->��{vԂCs�M�ƽе���7��W|{@�T�^a+:V�.���r9�@ULך���{��;!��X+I��FR��Ã=%�|��%�L6_դ��5�1A��e0�����{������^g���������]�^���0y%���A0J��7o��������f��5YύΤ�D�9���`e����e��i;�����0�C��	Hk&U:����Fѳ�����~��9eRE	�����Y�e��P>Y5���L���&��OC_�uq�x0�V����KC�ȩ ���~|��+�e����\1n�'gd:��}:���_�wv�)���o7% �S^A����,� ��
�§E�jy�|ױ�@i���Z&ac�'�x�ѷ*W��:�*W��$��q�����eA�^'���7��J�Ѕ�'�+wj\�C52T-�xm�	qt��8�rR��5����]�µ��,u<o�̑h�H�Q?���'bE��[z1����}ĆE�C�)X�Ch�{c6�}ine{k�V�=��1�Vn1ahb�w�☣B�t����l��I�k1�]H���BxiN\5�Ca�/��)Q]��_z��L�e:�x��9eqn7�ƹ6!�A%+��fI,5��8gʖ� `�F�.{t"��{���P�WZ�k�g�@�'a����K_����7��������)����|�E�ût9�n�.b��Z�#�܋$��;{t��BF�<&��-!�����k�,�wN���w�|�)�N �N���>���Wº2����ei�s�}.��!5s��c����=��
)��,�����a~+���m����ID�j+��$�,t	~��%�\�4}��]m����Ri�W�����	��w����F�$�펤<�8S8�N��<q�1�[��5c��o#�]�[�� ���v?Y_�r�~�+lԢ�0�%Pym�]���j�yu��V���A�y�F�W��^���PzS��<rW��dlp�����@�"z���ǣ�u�b:���O���ƣ#�~��*���r�����ߨ�/���.C#U���F*Ű���VN�gҹ���|���>����h�?��z��O�[M���HKrժ�J����WkF?<��v��e�I{���'��FO����.��$�7+Ҳ�\Z�yo�P���C�A���+���,�}� .�i����k���8�,1�Fa��q�iu{w��X�D�ڛ����LW�v��)O��˼�$��bך�_%%�������y��ҟ����[��ӾZ7�-�'SX'=�����U(��9�\�LTĶ������՛I��^�D?(�@jEq�E��,(>Iz�
V�*�y��W͔�v� ���v_T¶�#��`~����������S(�Zmǖ�����I7�:����UR�S&��)�������}&����,=�{����dqP����݋���KL-ӏ�ĝ`6�����+���:�"�h+D�3����E�2BnWv���NKz��ݥ�[�M8i�B�ג��4���G�3F��xd�V*��10�U�=������Y��H��o
p�'��E��L��ɏ%��qF�1�fj�WԔ�Q�;\p���2�?1\�"������q�8˕�����3�`T��b�*3[c��5��R���a��(���U}���]�M��#�]5||l^�nV���u��'l�Q����h�O�'����J���o �/��)$�-}���Ѽ�o_��k�~M��.�1�	]~�p<j�4��������)��#�9d��k|}yTLj�6���/�}ޏ��b��z�dS�1��;#�O\��A��[ N��e�� �Y�B-�(&	�y|���.5� �ca�p�|^V�� .~.�`��2�qn�9�T�_�Ŭ�R�,qBmJ�*�
��{cE�I�H�=ӿ�¨�ư��ݜ��{�Ҹ�{�Kg�u�#+�V�����9|)h9�J�!"�2R�o:GS�1��d�:�vX��W��eA�)���d�zu�Db��տ�X��A9���jJCN.�|ܙ<
��D���?��V�{w[�`R_�t�ZoGBx��	'�����\�n�m���]�T��%���7�<1����΁�E�?���r���;3����G����g�w|:�bS��O[�:��A�?�7X .�ŧwy�.��ה@]�YX�M��;�P���V?��:ː�{� �r���͈�ʃ�Խ�������⋶�&���_�o�o�&��>�(p�T�����݈��/���]k��y5�נZ��I�}��(�_Ĝ�60�0S�+�'�����ti)����%��z�M��E�f7��\�u�����kb��:�y��=q�b#�t?{o�<��z��U��4��+�u�Y�t�|�r�l̓c�wj|j|��o��D311�d�yZnb���t���j�H-4@ {���m�i�	���W�=0Ťd���R�����k�\�tf+Y"X[�1����uಎU㭋\Q|�����a�׿��]��S�M�#66^�2�P����b(���_w(��=�N�lb�}t����h��th�۫-J������8�فӆ˰���*����|H��";l?����f'{�v{�F���`�0�M/I�k�U�%ҝ ��Yt71Z� �D���B����������� =����`��e7X��Y�R�i��k�nx�!4̢�^�8�Ɵd�ȉ�w��Yf���]��Xߎ�T WIL,e�(N"\d.@��C2.2�;�Uy�=*��m�)��J�p��|^Q�"���D;�a&D��6��ɵVr��fN٢>�����ӝ��e0�P��o��u74̩!lrė;Y� �J=$s��;kϔ&3�x�碻�/ 8�/��P� �$�JPg���ey|^������%#R-�>�a+�JraL�Γ�d����|�fk���C�o�9T�t��B�	�c��R�W����!�,�͍����ԕ�ᓼ�Ѯ=��,-h=D5�>�>d��8��z���&1z��6D��4ݒN�='�?�&i������(3OW�/D{d��2�<�=��"�6���g ���7�(^?������:g�F����7��I�}&*/�4Xw����.�W���g0��3�%q��r�V��ڙY��r���˳;eQBo��S9^"
J���fY�����Ҝ�|��"^^���cBl�{8�Lट��k/%p���s�����xMkr�^��*�s!�Q�Ћ�iJ��Xv��wSui~������X"�@���W��was_���Ӕ)+�ؖ��9���vWN�=-f٨��|ɦ��$Z�^:"���o嶰��,���tX�����?������I��pwR��Ƒ�t��o���WE��!���3嘐K������^/�氬M#�
I��5-�ˤ���fa�P�%�q8?5��?����@��$$Ҟ�Y��o�aO��Ӟ!#�#���0�vʁ��w��V�:WٱbX�)����>~��]S�踹�^���L\�aH�����}�17�ɀz�V�-`�4do����^�f�Z�d˞��S"��!�˭��y}�*'�Q-7`�;�ONW����Z'�_�n�1��ho}J.�Y{̢y�(�t?���L��-�B��Jwk��z�-G���,lo%a�q����f������VE�R�$���m%�%�ϥ[/�vw��z���D"�+=��&Tۺ;��(��lJu��<�[�ć��=f�|z�Agm�j�m�)�E2�˃���8yϭd�'O]`�p�j�����p�.j��e��m�ظ�.��hL�;`�P/�yV�9�G�P<lf�G��0qN]�.'\��H^�)0A�)�)%�w��A���z�顑�)X�$z��7*a`xҟ��/�Q_5'X_�'7&+�c�dZ=]�f�.[��k�������见x��N��~���-K�7�I?���vb�!�/V�~H���\;6MD��� ��������ӳ�k��
�6-U;�5S]�҆.)���Iί���T�geKզ���〳o����b�*]y�>rJ�
;V����#�bz=o���	�1[�n�L�\z��waD����덤����%̵���Ew��O+�ew	�h'n<�C./ll��*�ϣ�Nj �oVϽ���$�^�j�W
��tL:���\w,�X	~7���	@(G�O��v�*/?�P�Dͥ��M�ݟd}u\�����~�Q��6L�bS�2Wn�&����P�;�jsp�S:3�&4cTa�Kaj����f��X%-�F:]dO�
 1ޔ  �^
9�j����w�ߛ���a��;+QP��*�A�+8��`���K|�āEK�!�nn�����}�����Ml��=jeߔ���\/�j~���4 ��q�|-]�d��Q̕����a	f������xm��ھҟ{��L�NܟVB��ޝ;����F�e�"��n�ʜ��Iq��ݭ��ܩ{��#�ŕP�L-��	K�M\�⽗'��wo��-����d��c���m�L�{�<Aߏb���˝JRz��ćW��V#l���ؗ}цN%L���Ɇ,i�!�����ꝕ<hAϸ��sU� .a�j�	�`tW�%qp���J�F�ݍ4� `�t ��/�������G�/��nlW��:���>�i�b�9%t����_L�Y�LaW��Jx�Ö0&5�P��I_�7P ��D�:v-����V~K��۴�W͌a�z�c|��V�Ѿ���9)�\ش� 	�3*��bd�(����(�by��f�AD{��m{«#��E�l�C�~`������읥�29�r�1�B��cØap����r��/�ȏ�0��j���}m�mU�\q��=�+��#[U��8LP�gr*�ǟ*&�i-�9��
\�<Z�O��;��B�|.�.xuL��mn���g��P�s�l����|�uzh��
I��,�чn��%/��u��~!V���R�$����S_q���V�Զ���"��\�9���w�r�����j޸��+?|��#�4Nko������@��r+6��:�{��a�K��i�- �(�/`��O7���e�{��/�>Ӽ~�l$��1��4
�t;JѼS��o��ȳ���d>c�N�`s����?���YL$g,�m�^g�3�je՗�o�>{����L�Oֿ�]G|�'�-���	p�i�4���
1���D��pjUiB��TլU �H���e�P���kԢ*c�%�,K;��	/��_̗���ٱ�B?�����@����0�Q�`��=�Bu����٧��V��W<f�lp}ny�x[���wa\�=9u����,�͒�q���N?kD���,�$���ό�;�8|c��	aᛴq�x�ȫ���Wt����U�e�`��x��@B'���
Ӥ�_H��^Gݬ,�B˥:ya��|u����[VNh��ڼ@��:�S��tq$����3�诌O��^|��)`�Wh9�RP��ϒ,�{�~Q���Wg�}S�����B߲������Tq�I*+h��c{�y|$��2r+y8'z�"����*��L�4��"�ۙ�E��Rm}v�4�K�k'��C���)r;�X�K�x�]�ڽAW�a�+��ƽ \d�L��d�k�^�=q�����k%���>��B���זi�(�}o8����EAf�6�Py���5{�	W�<?^4
d��������ׇ�����G�E����C�Ɨi�T�eqZr<���^�ŝ���v)/b����3As5^��"�!�� {��ura�d���bD,���_A�g1ψV��Y��	�g������y�R@W#�?Uq��%����O� =N+Ln���-��r�	���o���X0YN����Z�qq��hy��F2c���U	�1���Д��U��P�㝏c�Z�
W�L�ٰVm���x󚝞�'x`�����j�G�O[n�s�3SU�����W�שqt�ٯ�9j��xz�Z4�	r����lN���|I�:���5���.�"����DBէ���)9�O��X*���b�7������qt}�sHC�L�͙`;��9|2k)U:�t���y܎�Nq��ץ�@��@�7o�W|�x���L���Xx�_�\���Zo�G���nt,��J���G�QJ���"}p\	�gGO�,	�K\�f!�D
��� �V��ɲx�S���o�����{�[��k�)���*���+� qc�Z�0�+��<hO�c�/�G�q����W�����S�=[�w�G��v��D�͋'{0�2:B�n�[���#�=�P��'�0�P²�i0I�
J��C0�����鵯}�#�I�C�<?�F����w�i�l���:����i�r�]l���E�ù�Q%�b�.|O9��ߦ�� y&�dmf:���b�d��=6 ����`<n1JP�[V����YZE�#c����p�#�sŠGU���ˏ�BE��a�u����h5e�L�*�(�\��({��_E�v�z�=<��_�,�ߩ�H3FG,�����01�P�3�8����h6X3�+�%G n:4�����:���2��bOP��4�|I�
��t:�r"�V9)���(D�\��ةv������U�����ߘ��N��3ߑ��E��� A��#�t��v�� ���Ga;��)[������9�m}(N�8���j�S��W��;����f2y��(�[EE�K�����K65�d�ԾX����߼�s$�e��f.���˥����Z�,"�C2��s��eY��@?�K�
� +0�Z'�j9ss�6��V��t�/�~Y����h���F��b"v��2�97&��d�o�p��C���ӡ��X3��	�|�ة����ϧ�)x�[0��b-�^�>~��ļ{k��k�Dv�ރ���%S��Ҁ�wKi���g3/�^|[��V��|(�al2<����p�^c��y�`����
i�a6$SD|��Lq�m����G}c�)$AT���P�یT�b����_?Q�UC��pE?|�6��Hw����e�[�&��݂�I���6��~�  �݌���ǆ�%`w�2���hCG�VSL�S�oc�th-6u8���=�/����0��Hb`$yQ�CC�~�W��ڵ��Nk���/x{��}7!p�P�i�w��#�t�V� �� f^6�v΄qE��ڙ��zsF����Ý,��J��#'��ԈW�E �ݜ>�dȗt��<W!.�n�)_gX�(��B���dW�Yb�|���K%����z����e?�I�r\{�Um$����(�̞n �s��jy��"f���mT�'�Ji<�#���4ʖ�z5��*�^X38`Bi b*�-���"·���]��UC�ˬ9
��<��-�D0�y�R����or�3�I���
Q�ͩ&���1�"��؅�*����n�?U�2Z�"�w">�՛�{DM#�Uf��BRW�������9��4��R_s�*��L?�(�w̾-��8�JX�Ƨ�#��z�T�뀛PД�I�Yؼ�_HK�R"�GeZ"߰ �w�@ܥX'��r8��j)Ki�O�P���' �C��L&K����w��={̳@H!�%�5�m��o[ę� ѱ��,�l�ƨ��� �L��\7t�&�֣=/Ͷ7o�z�*A�I'�jLA���3���U�+����i���Ȅ���[|�����q�l"�t1qO�S^ X%L��t'͵�Q�)9�B�j�v4X�m\�� ���=h����- .p;�{[�+  ?呭��@g���H��g=ҍE��;=qA�6����#�>r#��:Bg8�~�[>��;ˣ�M	�3km����#Iߞ^��Y���JmiG�!�P�c ���=�8^�B��W>3�".S,Q>�y���ӵ{WϦ�V,"��2EFF���O�RJ:d���O�^y�6�Gn�&w&��di��X��N ����1[|`~�|�~`b��a-�eB�� ��p�	�Qo�':�'�L# f��ȂKa��`��7>�����^EL���xxi�޺KK���Z�}����k�+͍��gcv���/0Щ3�޽yU��SrV����OT�X�_0E�rr]�tKe蔛!���KT�c���ϗ�S��=.�c|�<���S4�ߍ��9��L�4���b����.(����E��|9T @��:���3p�q1 m1EE�l˥V��0Qp�������������K�_�˯m�LȐ+��.4&44��L�r}�͌kG�xI1�;���6�|Wr9Q������t�Z���6���l*���XO��-_��n����~1���ը޻+����E����4oܮ�a��o!����P�_�����d|�i���LS���r�8�Ը��+~��i�d~]bҔ�����ӧ���
b(�K9.����J1 \��F��_8?ar��]�O�P��(����}�0�X�� �:{*9t�#n��Řh~����==:�p����.�0� 4�>�*5a�_ےޏ��DSܹ?ҧ��c�g<������ivŽU��T�`��s��6
�t�72�<U�`w��%�Hs��ܽ�6j[L:���FCz�����V�A�
��XL�u���67tåRVo��N]e8��?�UT����Q��VT�^ȁ3�f|���(�EM�(yc��.U|\b��AT�W~���|�!��S� 3?.�N�h���#�z�M���?��%r��J�4�M~j��6�p=:��bdVlB����Qm� �E�w���Hx�o�ʞ��C��X�1�?[���+��/�Y
"���$�=?�#�E�3J6�f�J�X��ꓗ�U��
6�Эm��u�!���Xg��-�U�^����pw���h�φ�wh�k�P]�Н�wßWt;��&��Y����5c=#?`��V��ν J§�6�5�/�V�ӿR�_|�;A�A�� "%%]���F&AJM?� �:]����[�>��|E���H�;Ð*��Ť��e��U���5#A���o��ݔ����$��^������ j�@^�q���48g�F_�H_�`��g�=@�X�3��M|�����j��B���g�gZ���}�;�\d���-������
�r\�n��K��V����	mm�z#���aǬ��$S����{���^�@��s�[�PUd�t��D��N_1"��nA�ȸ�nэ�*�p��ՙ[AƯ�C�xx!���	K�/���$�:*����M�7��4�Sl\�W�ҿ3mo�&�>e�jX�&=�͕��ܜCT���+t�/��]�N/�P*���<�>�R�I�1�!�S����'�����-��a�h�߫�Lu�>���~�J�?A�'C�[�E@Z���Ȏ�Ϯ^�Dϸ��	Zl�f~���V��L4��� ����\u��'�h�E&$����E�䫍�oM��?�e���F�6�қ�{�Ҏ�����i��MH?w����}JY��W��B���I����n��7�0{Μ"{��~㎾o�]t�?�+��Iȕ����>��D��<W�$��	��A\\`�naAϸ���Oƣ�
[�� N]>x4�k.�J]��:?	jٵD((���2�[ݵ�B���v�`^�ՊbiôI镙���r�`N�R���������x����N�1Z�q_"6L�������5Z�F��f�v�ɵ��z]ѫ%6��]`){���IJ���03�{*����`�y��k�0b�p n�1B@D�";bd�����&Mj���ퟴ��)���w9y�F[2�Ƀ���`S�Fq��"�a~�����$CPBB���<p1=��oF)Ar̯H5� ���zvN;�(��s�����{��eN��z]�@��vv�*�ۇ����fj0�{�Q)r4��Uf�L��e>h����0B�(���	�۝!��8W�����]�~H\����U�����5�R+���ڂj��?Dq� 4��Sz��᫽�#�Ã�|�	��.K� �s�pW�iQ�K+Ťy� ��q�7�F �6I�w���p7S���n�-���#�B>e���ou�]]�j�L��_4W�������b0G�"��3|����Al-ܖo�zt����3�eֈ43\f��e���S!����[	�*���o���\�����{��`�n0�i^��|T<l�D4�%�G��om-���L?�����k���������޳ۜ�u���g�]�ϽPJN�)Wu7(��b"Ri��Yf�� ��(C��}LM�����.�'z$�`���hLF��dA��Ð���,�jG?V �F*�N�@���o0b&�iW��k��9?Z;w'���w���}�Fm]S���v!���/��}c����_`�˸|�2�fv��?g#nk�bҞ��I}�Of7_�q�� ���bs����C�����������8�Z\�t5Z`��:�E�~t�Z`��88��z�f�A��e>D]`"�ޑ�#maGu�U�o%����'),�c���K$��b��-�N�oYYS`�J%�όF%�e�0Ŏy���D��گN��wݘQ�J��)�����m�NM$��S����ԗ�C����TdM��B�d����%�1�2c%K�ױ*��L� "�0c�nB�i,��������}��1���{�s�y����y-�be�܇����`��eZ�.�qhz�C����h>��c��=�������a�9�3�c|����=[�ȋW��p�$��8{��b�6
Mr�K]�>>��7G�������_ܯ%�}qZ�HkW��2W��v%p\M��4�p;V��҆jbʆR�v敘�J�k�
%�}�@h�(V���l�K�kc.L����,�� L���Us�ҷB�	9zUd�~7�G��|I�`��"�MLRp5ֲIW� V��U	��d�p���"����:xِD�i�˦�J�|��,�$���=M��'h�.���e.����!<q�Y����֏��w�S�H���bPc`�֌{ 4bP}�r\�H�~y�;w��K���ㇺ��'x-G,�Q_|�i:z�� l��~�V����$��"�s[ ��!����nY�|�0w:$�q{S�;�y+'�𧨝�8�l���,'���/M:Y �/J�{�2�c2��sT/s�U
LU��8�dD�mw��V�T����Ɉ)�x"���Q���'ܡ�:x���kY�����Z�&귱8Z��|�K�Zw�L�P��V��rZF2����z"�e��
s���[���B�}n��Sw�'� ��	���=���{��W�WX��8�@�{�C;�q��z�U-�\3Ӟ��V��#�)j:[��G$�3]���*��-]�)�k�0�k�W�����|���ϯ�n�ؕ�~Ѿ�C�ΌZ�J+A��x%��ΰ���Fϊ=�E^��v<lb��4���1�2�J�Sz�A��ՁI_�#t��f�5��%����Dű��4��!�ϊ[��DA1��Ā��4��a�F�_6���]�wH���*�Q�::�z��3[E�Ep��O�Q��b:� �G�^r�OǭY1��Á��P����.�[��<C�/8��|Π*��V�M2���3�qz4=�f�iz��.�h�ކ�1�kd4��Zˇ�.����i9h�^�Its"�F�཯e�N(�`�!�R�z���f���p��S��T
e��ü�� ��@�K�>�%ϝ�vA#��c��Z#�l(��;M|��ӟ����m��䄿��8�z���.D��~n��.�����L��O7�]l#��L2o�8{D�n��+�����Gu7=����a"���A�S��ޒ3������k���t�,��!Y!>f���d�kn[+D%h�~<���yfx]�xB���Q��U-�)�M,\�]-װd��*Q����o�����]aw�^ybʗ�=����a1�<������be��i�Y�}����e��c���#�þ�!W�~�0�~>��".
�~��n�V>����}XQѰ�>��8��X/�#�ݵAoWf��Z�����[�mOCV�C�Z�z{�w� ⌂�O6��wkY��(p���A�S��7ɏnDK�5��)ϻ؊�����?�GqW�`*o����l�s�;.��d������ͅ��V�Ч9�ɜ��\�!���i��Q18��@[�x�/�KXg��ԛ��ֿ��]aL�>.1���n��տ�e5��t�׃�םdVï~����ՋBgބ�)M�[���藣CPgH�8�����`H����+`�[�Z`��p$�*�IF�97�ǖ�S̞��
�uD^�U6k5 ��/߫S������ą??/,+��M�kn_����[��|[`����l�)��7���WDC��ɘX`xX�k��y�;�]t<R0�u���]F�]F�	uVІ��h?m �N�ӵ����lT�0�n����"�+��HV0T�`�_@�=2�?�3{(��B�j�ՠ�H�n(�a]=G�ZZ�������q��_:��N^�&��Q�\g����F���l�Ĥ}�Go1�6�����}@���vc0.��(u��¨cv�jg��%��d��I�ɲv� �]��EQM��;&&��u<�k�zi ��ٹ��Y8�Z$
P|J����0�~A\��幼��3��Vv�,��<	_1V:�ֽ�;��%^��6����y�aH���ظ)@Ѿ�x$��l�\�"X>=��;F,�`����^�[э�ٯs(
^���3�N�#]����I�w��F����8d6���]w��'i(��~$���+-'��'L1E'̵�I�F�K��s��E��+
��KY�	���<��oY��Z�3Rj�
�l�W7�,���[)2F܆�bG���&&�x��������b�dL��:��^\x�K��{�;���|$��H��P���1pک�a����shd=p��Ͽٝ�d�$w]�`.Qk�%��+&y6��B�\e~`)~�`��Yw7��ܸ��*MϹX�ggk�^hO��"�ܬo��Jౝ�}J}���4��T(I��f�g�q&U�K�_��8C�~���m�ZXf��_���J������湃�����~����o��l�)͑�1����`Դ��K,q�:����Y�t�p�{�փ�xp��e+��`�ފ%���y�]����Ѐ��>�z	{��>`�����^T��Y{z�|��,�e!�+��-.��<�=z:�ӭ����R0.�}�$��X�(��	q��-?i������\��쩜�Ř���]�<O�P5��{��� 8h�r�,^_��%�$�ou|�X�"�=�[��on��"�)[��ߋ_Em��=s�肖+��6��� ��(C���f��/�k��7�
~�s�w�h�d YP���o"$�����(�үݪ���,Yg=��c�(Z���Ih%�j���`B�Q�` S4�T��o�p<"��Y�
1& ���"g�x�K��
����%��Le���i}��8��{Γ���ɭ����z�{��4�LW�OS�Hй��0<����_��"cW7R�
�C���e]ꀴ��#e�ڧi�_]��uUh(� �)ul}"�?D��o��-0�B�+>��s޾ބA�d��d�R�}7)uM�ؙ�6��
��0pJ�U������S'����~ ���`��ޛ�ߚŪ4K�o�3����S/�ie�E���{�[�~ȇ���hǁK�z���<��#;?O���/Z����<CU4�A%D��4`��__�S���(ʚ�����9�-��F�&af�����ĩ��� �T�_��s�<��}��P"Q��k���˸.��i��N����+B�8�7�eud�����5'�y�eW^��QSC�
I~Pf��܄ӎ��,V��O��e��.�n����}~$�|�!iS����!y@���qJ�EӃ��mo��I��%^���1b8�H.��8�"�n�=��E���Fl�_���Q�5�{;*~#S��O�p���%!Hk׽&K�׳��>� -�77A���Ԥ.�]��%C�؜L�hXE ���S�M%��+�hB̈́S�w&���T�MԜK��6+R�8��1�s�~�pl��9U����O��� ��^�cix�L	�3�8�@|�M�E�/���~ħe	GT��9A�S��[K��W��S?w�k���H4�T�lp{,y��A]���'�O�P�lmt>h.ӵ"���4�nm�1h��4Įq�Cn���CƆ���+�y!` T1\ z��,��Z`��8u�Kio�JÛ$�I��~�P�a��^t/���ڇ���\���$�s��@�������	U���H��T�;O`�� U��=��y�D��G�:;5��q��5��W�3X`�w��]m�m �5ܣ��FD(2��BI^.���Y ΅_�B
���fh����@�eXG�G����d`C ��C �#�<ݥ9*�
��w$��J��CY�eB��C��-LX�	���p��T9I'?dА��k�H���1����.�`.�f�dz�<�|�p	�&�K��SS��_�P��u��f��x�}NG�|�s�g�l6�T�	�
�;t��ٴ�����[��X��2�����UD����H�M���1܂�o�N��(�,��'��h���f�L��Jo��M~��C���'��#���2f
DRƛ�GZ��K}|S��k&D�o�� 鈍�O�m-� ��늗��H%�/�9?`Bp'��f��",�����k�JJ�2�. T��A��S�בK�c�GH��֍r�h��n��j�����:�(��/�
1��o��nY�?�p��aL�-��l0!��� c��G'��[R}n�&L�7����ՙ��˵5���4����N��F��F����D���
��K����n
hZ�-����Ҿ�;���'��(V�����	ᴴ$��·�0rYΥ���������xT=��`JK�s�6π	Ҩ����S�`y��U��~Ϯn803�=�Z#w:_���B?0Ŀ�����b�~��?ׯ'�|K�5��#q�Q��3φ�jV#�-�}�l�wc6�7=�Mp�.ڿ��U匿0��$���o�5�>����3�S=k��tH@-?�mV��>�(�aҍ�>E����ȅ��)��T)N���y̌<�s���k���s���[��3�W'O�̉�-��_-3��{�K� %��"�\��u�
�H�Y_�gk�!PV�/��h�tn�cТ� ��vq���E��?��k����� +֤��ȁy��2q�p��^w�<��+�l��ݿJ���E�=�Խ	��~@�N+�D����%PZ��qǩv�J<�
Y��K ���c��>	P#�)�E6
�7�e�����u.��8�Y�y�.�$5�/�c�c��&3�q__�����r���f+|�����	) �̻ �!yQ�P�uJ� :J��t�{��A����[ھ�uϋ%	ʘ2�薖�����[�
�e�/T�\�$�%=Y�(=f=�"Q�h��D���(�e�o��D��8~�E�0Y��B�B�� ����0\�v�*vW_��
��M�CO���e���d��8�C��1ϥk�Wh�b@�m����Ҥ��Q5���HqMѮ3��"����dl���L�lH[�0��{��>��+S�&H���4��������::סu��wy��B"��E��$�LO�{���\Y���`��Cv�ͅ�GJ�< :V�0�ϗ�J7>E���N�b'�}(J��7�+q��BϝvM�I�0�˦{8=Ε��gNe��n3V�70k�ZJ�v���E1���R��Mxͷ��u������፪��ͪC��S�&����i�i'������J��w#X���r]��Z����mj��(��[5C��F��,,���ě?��#��_x��G��ȣG�B��̗D���z �K��� m���2Y��w�Q>�1�Fd�����R������5��~+����ӰMK6+�3?>-v���VsՊ ����rU���(�y���3�O�g|5=��w���woc�]��)��D
S#w[���tMnő�n�ř��$�f��=�m�J%�b�ދ\���ߜ�ߺd�S�����0"�ؿ�D�)�������:~�{������{L*�
uZݐ�p�e��|�(�/�]��r�	Y�W��{���߀vYN�%i�J��^@/�	�C�VثĦN��d��z�_4g��&KG���lw�c� ��R�m��M�T�I�����)��{��A[�����7'�klZy�V1$�:Mhs�G�?���"��f�ы��Os��&p�
�$v�B�����#���������O4z�elL��yiҩ��h5IA�Ρy��=�I�K$������:�;�u��3e_Q�d!DS3k?�	.���t
YP�0�M���B�0:�"�fQ���=�M��W��Ʊm��Mui���A��S�K�3���A���o_0Ԕ����|�����/��f�	x�tP�w�ݢ[mB���v��
�o?�{��2.3xv������l���]���y庬g�ھ�����������S���+�b����
�p��Ý)�����-0~�1{6Y��w�))���
&����D@�����)#��0o���	�R�\%��W	���A�pš,�䖔�Cк�th4a�Z.�ў����,�f�w��վ�}G����G]U�U��p�+�|y�#<�<,H�w�`��9�����m0V�7��}�S�p���l`�T�l��)����H竲�֡������9vg���ּ�?n��U?����q  ^U��-�8m��O�(�b��^�t�p/g��I:T�s�2H��U� ���;NӖ��o/�aG�Y�W� �ќސ�}��[� eͿ�l���G��tĻ�Oak��s���"Z���4�f����՚��
����X��8����{(Q�^��/�k���b�s��P�Ҽ9^��
�R)��Ҫ��D#v��7�s����Ic���&@rl ��iW�:�X+���$Nh�Ŀ��F
�S%B����)��B�V��]d��᩶T�>em�AwA;�F7��ã�q�ѩng��H$����o%zQ��э�>
$+�;�U����lȑ���(t;��j-G�2&�}���7f�'�����<��L�����
J��9 [�^�*���'h͖a��xr[��-M�Fڄ>mE���%s
{��6~|[�����uIb�΅���aW���x�k�q>�?q��<���M�4��
ӧ_
X�+@Ó�l�gr~�t<�(�׸��S����\���t�J���:ݾ��V��������mĳ�9�K����$�8F_i��-i�����,ۿ��F��ΪD�|�9>ݬ�P�Rp[�
`� g�=&�E���W,P�d�+s���'x���S�L����
�?�a�)?Rf�����a���C�*��w��Jp�I���9�x��3�L�2��F�����	����`��Ru+� M����DixT>�����E^�׬�P�����}����ZM�z�K+MO_XS��_"o�+���O��a�Կ�~���6�0�jނ���`���W���o&��,E���ͅ
n���%X�` ��E�l�,��}�*�>��Mg3���3M�i�J\y�W��&�7�F� �%q1F��?����@ӹ��&�	��qnqᔌ���Ǖ]�w$lU/���-f��(���no��H�w�K���cgsD�T�\�(a8-���c��V~����]Zj��E�`�n3��tQ���ᣏ��p�'S.��E�댛��.V�^���v�\�F��������u��*L��M�gf#G �#x����xו�)�}�:�N��������2+c?l�ε��U��;]K6ʮ7��)���~�L"x&_��HR��3���/Z���7�]�����%�}R��[9O��K����TV�w��7�������䧟A��J���p����������2fI/�Ѫjɺt$6�ʽ�a!�| nj��xҼ�ڃP������/ c��P��g
\��,��J�|�5w���t�bo����*���q����:�Ѩ��H�D�U�.�6_�vJ��-��ə�L����۫��̾�񔵏�s��n���Oeq�Ϛh,�N(��ܜ��s[n4��gΚ�����E\T��fR��፿���>]�f���g�|��h����^1r�9 6kr�h*����Ԁ_;��9#�Z�+��eMM�rSEwi�0�������2Ȗe����̍�`�%�;��°n��p m����6�~�7�.���݋�Z��y�EU�h�z2�0�tp����ܷ�˄�l����d�XO:�G �G`l�Ds��YM�N����mV����fAH}���q�?-kx6:ӳ$��w�qg%R�sO�Ω�JX&i^v➸�Y�U�������d�?,G{��oX.F��g|��K{j�fFq�=��G�v��p	.���|a�����S�߿Ij*9e\9�v�_�6ω��|x�]�䂒}���ЪDЗ<0�e�����U��9!���I�r� xF�TT�?�]k׉V������L��aVLw��#��L���	-�cc��0�]�o�²���Я�R�o�<&B�Y��_��u���h'W��~��*�<�=�KBy]:��bEɭ/q5
tp��@^3SB��U�,<Y��a�/-�74h�z��҃{y�U I�6�e��iX���#W��F���e��������Дjf���4�W�={{�e���F�\y�������l��6ܵ�+Z�w;�KH�}~K ��tvMYP���o.Y���E���l��;j�'K�쥛�A/?��@77�ş��E���G�u�g$b�fѦ6��}����v2:͜����#�G��T��;��#k�_(�X�y~�!��=g�z�z@�4塀�U~�β1(�bɭ]Z��n��c���PS��$��wv5�-�`�٨k��K<x�(����V���d�Ѧ�4rb��'צ��N�=�<	���Y�V���P���m���o{ ����k ���c��t�qͭ���m%���W9b�?x7����q� ��h ��3#��˲�w��S`*�e])��*7�33O���[�| S �m/�|P�tT�{�0�_�$�?�����5>*y���
g�Պe-g����.{	�p�;BO���P�oXR*�lt�Y�XhT&��}�[�����|�Oޡ�y�"�h�J�*�E���T�u���"ZU�Y������G���Є�~�g�1��{�Јxs!>T�C���~ܴ@�8}�}I��X�!+X+~�����As�� �ڔ�������u��bG�S�ޒ����P�F����Vcje�#Z]���C���k����ǡCA�Ņ�Td��0 /1�Aڠ}�u�o2�����GK�2��ׇM���T�j�G��f���P�)O�x;�?:G������6GA(Vb�X��-��v|��`�+�/��Ε�d�,T�����?<�9�L+x��Wdؖ�/��o>\���:D��F�1����?'Ev]#�m�	}#�ܜ����x�V�yz[�|`�^ ����b�������E�ߜ� �BVg��i� �^�+KD���f���O�s�ٷw��J|E�ڰd=O�t־��W����Eqϻc�f�_a*{6Y�Z�'cK��ӏ�Lu~�6��#?���"�������x48J������#x�٫�Ԩ;etT���^T�BA�	�����ME$�f�5�QPN�,w�^��P��C�D��u%��-��v���p=��T1����r��(�}$�r9���D��W�K�'H������?��(t���p:�1��6��@�F��t���ޛ �5AK*�-��1a~~��>���V�m�Is���?�߷[]a�Wf��Yv�{�
�Z�`��������U}��p�gYc��*Ӭ�	&Mq�I�4.����tTL�A����ff��"�j�XN0�y�?��l�����#��������oG�8���睒l">�6{���{��������J��fb�\��o�w�z$��	Y��z���M�j5ƿQ�oFxQPR��ҒH��~�[{�����m���cL0(,�����
{8Kb�U�ݲۼn��i���I\ƶ�y���:\.����]AG�~E�� �/�6^ꢾ7�jI\��xr�w��k ����\%MKG�υY��$�82�Q{+tNZ?+3]#b\j�>g��{�3`��~W4�����~�2ʾ]�~������������Q`�H��I�`���Ek,�ݾ��I=x���X���~a�6�E�F�ky[a�[��+&�E+���� �_�81&
����v�h�DcD��>�B�v=�+w��DJ��ӻU����W��b����d�,�������Cd�T�	�D��g�FPL�wM���&Lez��.i-A�:]�̻��!$b��|Ii�{���鬗X����q7G�����<�gN��b����~�=���S��V��s���֎�z~����`&���'��T��?�p�� 7 U�o�u����/-�VY�4	�|f8>���Ѕl��m��QZ�X�]��ٯ^j�Vp����`1ZF�N7$�3-�;��r��f��W�'���������σ��� �V=��$��pu9A�L0�Xۇ���:.�x����)�N�z�I\+���ݯ�����c���[c�EQY᥮���wA����pQ�.�2���_��D���O=bɐ Rc�Z��,�h����z��Ň���SӀw
�UM̳�,���x��_���b�7���#�ʬ���A���~*Ǽ:�ĝ}�`��)}�k� 2)������x��l4k-a} ���H%��� �����8#܎�����>4�%�N�y�� �,#ګD���X�W���F����~>�`����瘧������݁ ��XMV3`&�
e���KKHH|�ic�~�yN��x�1]*�Xp�(�c�%�۳���X��V��!T[�l������8Sш+��W������G �-�I҇eχ���m�yC�#�J�\��L9����}F��AN���X4��E�&�Q�R�hy�K�ܖ��ڥ��t*�;.��� kM�>��(`س��ϾZ���|��}A�0t�~!��=
�>v�Q���I�"=�9�n��j�5��P���A�~{�2i�����תz�m�� �}��"���>>����Z��mhx���E���r��)P�/$�r���!��ˇ�����lh@����L�֫f���Z�Fs�� �8���l����j����f>�PO����W_#B Q�U8��k�\u[�jxQ��vc�_�T؂?���I�[]@����Xb������bx�?F�G��T���B'����U$��(\O�9b��j�
=%��������blb�%P��eF��}��"�$�5+��'��5I�yM?|�x�3Q�&(��=�w�I�ʻ�2'e-��*�>/����P7�8+u���7,唦���Oc��t���g�c9ki���g���['ɢډ�xs�	;2R4xO.Wy�>�)�)[��$���YwH8+�=��G�;�OhCS֨�Js�5���k�Z�S�e��}5��bn�r�Q�3?��m�N�c'���,�4��M�Dt����&�D?��i�-NͅF��� �Ō4 n�AM-���G{Y/����<��+j��P��pq�ޅ�Qn��d�t��YR��?�R�+�}�-���8&�T��]r+��]0Wx����Ǔэ^ح"x�"�oQ/�oو+wc��_�'���~Pl����2K����@��ؙ��f�T�q��[���w�G��y=%�����p���_*r��N�0lSln}t���nqc�v�^8I;h�&hp�80���v�h㍿5a^3�-{����^z��� RN�'3��L�DD�����WPj^���u�R˽{#I�^RG~�_;bV.�.OU�;*N�1ؠ�	�����D!o+{��|���IzZ&g�9�v
t\a���R��/p®0.�7�u{���sn"6-�����x�x��X�~2��S&���7�X�X�	�t���M]T���;���Д��t�����#����ٖ�v�&���F�κ�`�{J���(�pV�p�v��"yƃ�����-D����`:Ë��q���W��e� i�Ep����e���ʱZ���������0Ԉ�,L��!�1���h���uMA8��}�-�i/�Sd��$��̌`��k�ޮ�v�"&�g"���GHƯ�{-uU�CsO�}4\�ζO[{	�(E��z���Ѿ���G��(
��7���]�e��zX��~4#z>hCu�v��FLK�K����R�^��H���e�k�7�<nz�Z�"�IՆ�9���_��N��_���D8�~?�"�z,0���h)��^_��YI�����g��07LQFR�(�D;���8 )�4q�y�t�w��QyA z�C|CQ�=˞͡i���v&^?�x����˸��?�t˽B�v��ƾp5�t�px0C��qp����]$\�W�����o�V������YډX��k�V�Zf�����o��<�l�Ѕf�Wi�O�
��BNPaBp�Pi������m��$���Y���l�-�c���6^gji�`Ƭy7~=�N�$�+d1~���O��A�.Zr%v�N��9����o��Ú]���_���	c)���LYd�=\B���U��)٧ɢĦM<t���p���y.�%�;����'�Xt:J��`0��Z�k��x͌��H$5fB�B��]���s��w�455-!9���{����:6�_������|x��ޮ� q��O6�� <���P���,w\³�Is��m&�ol�W�'z����-���o�ܻ���;l�9φ #@�U�#:���_����_���B�ѭ����	c(<����{���耠1�Y��ӧ�:������l�����)��ls$�t���wo��q�Z^^~�?F(r�{���@$�<�'�r��j�^+�~�]:�논(ç|Nn���n��������Ǚs	��P+ �C��i�p��qn��+�r�=�+I{2���%�f�`�­�-1��_��#�kbN���Z��+ˣ�	��5��G��;��/G�&Ђ}Ч3,m�-t9�����=�Z�d��h�u��\�8}[0��8<P�B.m3G�3��5L'����- ����p53��V�UW�b�K�6�����
4��F����.7 �Tml�*>j�}��ZY�z� �r�F{W]�t��әѝn��_��|����÷�}ss�$�<}�o�ZG�?5ީ��/i�R0�5���"A���QPL�?\ָ!x4/�ΰ�S?NN���3���4�6�@��޷C��E���Z�*C��k��a���V~�vY�L�ӿ�ps-���:`�B��� ��oHs0�˼�Z���/�w={kY����d*���`���]R��2*�V�>A>�ݠ��͗7�l!@�R���K�$"����k^�u�K 3M�@9����0H�~>#��������g�����i������}����	�</�7����J�7�'w��_�CK�^nϤ%<�����������A	��?֘,��,QVkP�Y$��=�ϓ��������ߘ-�����/�< <�z\�����&�Z�m�Vw�o�k�D�aK@D2�?Y.�k�M�W�;�;�ѬǛZ�Ѵ��@�Ԥ���B�Ⰽ4���L\�J�"��㡲�.؟��b�d��8R�������e'��vsx���G5ͥA]���gG�����P�cx�})�u~��U��<��#C��_^c�<�_T���+8�.;*�����rKe荎y�G=��~"�{�Q���H.v<�"�0M�H��-L���d$k���X�9�i�[��O4�ج'����٪�˱�:E�.v�]�o�
�d[\X�^�����U�ƃ9޿s��%jhL^���E�U�t|��2�\-�Ju
R�E�9dcrr��"?�	�<ſ �R�2Q�LM�z��6Y(�׎�D�)@�AoO%S$Y.W� Fu[�bK�b��+�Q���@Cu��y�goo�ȇ=c�YZ���̲�J
�з'���)��M���W�I7"'��<<��*t9EN��������Nت�
���(�4�1v���WW��)¥~��RPK�Rk�I֧뙝��(z�����4�C�5$h'ީ����@�ߧ`b�+LKG=M�ߪ���V�'(�w7��܀�}P���Q��%e�D��I��6�C��h�|��4W��.�,�1)�V@�p���zԒs�z��(&�M3Q�i��	^PPp��h�i���(��l9Zƙ !��"�.�w����)����;.5O�y�6y��������L�h�qg��7�ϻ���?��_X�k[k�َj۟{y;�B�C��H:B�t$$+��Y�#^����d�{G'�d@@�� hB�h�\\,�Z�V�?s�ȴ�B�Ј<֍�0��i$�>P[�r���ϐR� F#2�d�u]
&֭r��"6�k(G2(<�:�2����R��[^j��?�q*��z�}Q2�F�¶RΖ�l�m�rU�g��Δ�s@|��i�$C2��/?'���˼}|��V��?�x@P��}>��H�M�
�%����Y%ۦ�$l`�L[ĔN��j�o�~�GGz��o1���%���>m�C都�r�q��E\�T��"�/ߢ�?[�Z^K������/�A@��W�*u��6�֝z���F�W�/H�j���l -����0��������v��4�^/�*s��Р�RΌ�(l7��u��R�@�E*�R�#CD5|ɶR���H~�ZZ-���ԉˤ瞞'�2Fs��+M�5b���ϖV�R��P<Z)j5��7���j'g��/1J�#�����9���Z��Ѹ���F����y��hU�|�|7�"DA�M~t>
|�1!$���}����-�HeM��&fVt��#�y|&�u�
~.����&턪#�L;Q$?��$�$��u�饅���u��!h��S�f_1�y�z�8d����h�<}{#E���|�8���:Pn	�0�1x�K�E�=o�۸�{l��Z�GH���U�\!�T��Qa<XI����)+:OZ�`�@�<ws���/&k�sOm���ᕴ~����
{Gb�Abuaaa�r�
���JJ)kGc�CX�Ud�LI0�˟���A��v�c{����'����ܡ�}�����(ǀ���kpr������ynr,dl�k1J�*
�()F�X���ʜ)k�㏘�O�4sof{֣�*۾�D�}��ѵ՟	����|�SR,��p��6𛐃�Xh�5f"t­@�#Q���q�	�O
�j�S(%3�ލ��W�����'(��.yyJX7�M�zl��}���ߟ���o�� X�`�Bι����Ec��LPJ���Z
T����*���K��e��򦮹z�m|�lo"Q`Bz�s�K��n�F*�|�)��G�h��
��:~r�E˲I�?�\[�ޏ���<��Pj����#b�7����~/�r�i���K�NW�_r�C$��]k3�C�H?������0�m�����m><h�L�nU��67C�	'�BRO�\j-U^�9��({^f׼��pт���y�VO�5m�D꒑��[j0š�m��t�2Q��` ��@��&2d>ڀ]m���������O�h؊��E�Yl� �p��),�޹)�j@GW��9*C��ۂ�'<�5]pÉX�w������JGX��v��@]��$���p�;1ĲM\����� M_�F��g��w3NW��Ʒb�'��DQ��70@���D�Q�T�c��^��ݜ�
a{��q�
8����i�c��E���ⱒ�xS�����`"�k�M�����^��P��JM�K�T��@�]S,�ۛ���1A2�O�>�5O�i�?{��>}%�^�����.7���Yzۈ<�z͒�=���*t��us� �!�R2tF�X1h��(ʖz~c���b�ﲟh����#0�G���Keü��f)U�$>�(��ve��s]���_�覩��B�6�.��:�LQ�y�p2+)����4���PYn㈴�D�8���W�1�+L7<��\���b���grAVz�#�z�(��9��Jx�PVIv=n3�f�*Lr������ىEB*)�n���.�4���MSOg�	C���8IbV���e�����OV~R��{��Z6X��B��l�I�f~Z�f���oR��(:����O�ڱ�q����#<�]F�e�i+@,vTl�.��a*M*�M� >��!���hE���P�D,�b�j�lC�������Xy�Z�yK��HB������� �ˁx�!b�R���VbX#�����I�����ݪBg����}pl�&ܚ:ߋ.�)��Dx߿wk*��R3qKvC�E���l��&�TH��ohC��p��:��2�xr�ro1�f��qT���)�����<2�b;6�/w�v���ݯ}*ʝ�]|�b��bƯ�H4�s�Z��w�p��ynq���o[J�jiO��~kZz�eF�w�*���	�_6 {Q"HIv����0��i��?|xFލ�Nd
�h��$�73q���]wÄ�0V@>��MDE&}��M��(*��0>5u����xM�P�i�~��n-� ��zk	9��Nu<�{2�^��wm�qzz۰�9*F�z�����x��V����y�7*U�v�
�<��-�O�e��[d2��$^�K�	?]��>M�U
|R�Ym���P�F觃E���8堑�\��3�)�l��<q1�ʙ�W�A3���m �}7���o��w]����6�N��Ð+/�Ȓ�	���dƖ���Ig$�0�"��V��Fw�O3��B��9�^T?c�WX(�"`&�t@Է0��At�P�����?$���ZK��cU2
��HI��)ҫ�6pޯ��D��r�|	ha�;�{�o���$I���h�\�פ��?%���<97��M�9IÕƆ��er�o������[&�>�j"���n�j�\��Yx��_8��5�)�w�١(������X3wGT���S__gB��ɮ�.�jT�ج@���ܨ��H^��3w�[�ʇ7�����y[Q�h����O ��]�;�-AC[B�1d��Mv�ϸQ���������I��}�s91����4�f{ʞ�h]@���N�f�÷N����_�5y�Z�����q�b�+�_�L��I6�߶Ec�BkF�4��沶����)��X��Q��i�/@��{��V���Q�����3����Q��_aj��e�&�L�WaI��3p�϶$���'������T}�X	�F��wA�nC����XK,|��,(X�e�倇��iî{�Ⱥh-ˮ��dS@�C��+�4����Fo�(�(Ռ9�J=,l�5�|��,�ٲd�o��{�� 0�X�}��}���rbO�k�����|(#tS�;3��Kp���#�]%���n:<�����盈MV�V�Z�!焵뵀�%PJc	�$h030���V�����n /n��^q\�pe�*��:��`6k��m6�%L@?�O��e5@H҂BҰ�U��iPt;��^�wF��8�����F����mW��u��N��!j	�������@@\G�(��d�WȐ,�42�j����'O��D��Pu�>�te�\�$��Du�)�n����5��2���-`=,�7�|o������OA�����X��[oe���֍
Q*����Da�Ice1�d�4*-
7�mH�(Y��diȒbl�d$�i,Y��Be��\�}���<�\5�\��Y�y��y����xǷ��|f�2����*>]�����IE��8��֧����!�~��&I��H��1�=jY2M��Y}b_l�s/Xj��H/T����f��� >���`�3����T��Ћ��9�/9�x:�dm���=�_�b91���6to
 `���_6�G�ڮ$���������=*�fF��&��1Ļ�o�������jd�!��j?b\Ҫ��l N���DX�J�����3
�I�K��Z(C�N���R�e%v�ƢnF����?#ث$/Q?�Q1�ԥΑm���쁟|\�z�Vj9;~<X�>�MA�Y�������d��������Z4<����
�DN����d�0nR,ξY�Q.��z#@�_;�%�Y�e'�����b��T�\��)�n�u��.�Xk���ICDv�k�/���7������w�]���`A�s�uww緙p��v[s7����	��g�F2St��Z}<h�z�a5�����d�'� ��9��}�v[gk?��i"J�͈r��+.�s�0�^<��$0`�~���b)�
.ܸ��������E�}�U2�A3���+t#8�o?���
�T0�E�)ݤj��r��v����������a$�p��]M�˕�5�)>������cL�g�)=��N kS4����A1��E����>����{c�%c6i�exX
@h�ԓ��RP�}ю�b���uu���;���TK���y�^��0z?Vp;������־|v����H턉2���W���^\�~�g!�����/ˑ��5X�ղ�D-'C��	��#�� �H�©�~6W���N�^�_�z�f��b �,C��W�ش#$}��*B9��?-�bп&A;���/N�9��۷����Z,���Q�s/�\���w2���<-�E u��t�g�P�<���u��2/�B5��ݪ�O��@�G�vrEm^U�rvUO����
��nl��r�ǥ����fB������}�c�D����Ϳ��f�:������Y�T�%+5���������4#�'o��1:R1~���ˡ^b��М�߹;�1����_�侥�p�>�U��2ٖ0��Y)������(?ϙbG�_���
w�l�8�!��(���e�!8G}�p8���u��>0��m�T�k��O��X!�o}7%��n��h���W��N���p�(�Fͯ���xq|5آTmz�C�Y+Df�N���9��L�5�?�AG�T�9������~��+��gӟ+�L����S��^�1��5j�����!@�7�1�d��L�rY6F4��ty���a��U1ܷ;{�Z w��9�Ӣ�ճ�
�_E�$�����1�K]���5H-�<h�c!�d��D�<��_����3߀rg�L�a"��3ߙ�Ge�|NЀ?�\���f�d��Tda��!л�D��2��Z�� ��೉6���^˜e!�-^�8j���?��|�0�NTGZ�y�n˨��`�Ebg�鏜���l֑E�L�%���1��W��K���݀ii�H���MV��u��6��>��u�X8
}E�q']ȼ&\i�'��b��n޼�����h�Z�O�ɰ&�Q�h �]A.�+��
<���S�d�G�r��5Cs;�D�����*C��i@ %�n�d��C��/}��e�u5�@]�	�m	g(C�,�+j>m���0�
�tI����F�t�>�p���>�渝]���5�����B==JM�t-Q�\���TM�7�ꋌ:����QS���W�\�Z��y�s�w�R��m5��+���
%�;F1U�o[lr�pQ���g�=S���/ux�E��� <��xX������y*%�Jx>����q�okY�4L�+U���^z$���dϭ��=�u:��Y���2,���KR�gTft�W��Q�1��{���9�:js*#�ܷ�@9���q��Ly��|����Ľ<��eW�X������wl��R��F�j�a���~��MM~�+��Ļ���¢φ�������*tPNo��?;_#Ѫ����j���	�@S�aK��.+� )������-��vA���zք�~U����E	?��nf'��l�h�mr�LɆ��J�g,U�`��s�l� �y���W^=�g��o����F���6fę��>��S4�u>����+κ�h���)��ۊ�zм����tO.g&�`��R�P*V)��Mv/�-����9�.�0���D��<� �l"��%e6N@�4�$������Ԯ!J��Ĕ� �f��>ê5�6#����Qr�]�	��CM~o��<m�3�6�;A��*u����ӚXeM�A~��|���[�{�x�/��L.J&�l���h�]�,Ң�Z[E0[�.���o���=�E���bN�bd�;a)���zw�;|U��z���Hi�^��H(mEA�&;�;ʀ���0�~6nnQ��+���ej�x͵���r��Ȭ���ǢE���8��ռ)A�R�vmdm����j�Xx[$:!]ȳ,��E�s��AY8I.[Z�<�Nkf�e8SA�	k~�F�S�p)XaRᚡzC�}!!�rUs�����E�����K%���\Ů�.��Aj8#����9%q[dy"�&�+?:n�w�F騳��� B�Ą����.�d���*'���KtS�&�q!(�i���V���u�� 11s�:G���ƥ�/Q=8Or欁�M�Z�CW��P�UමF��c̥p'_�'��;/μ�鼋
�Qԩ�t�{be���u�tF���:�Ih��Fo�2�V_S��d��fff�w.&�=�b�z�J�*U�L�@K�Ǣ��g]���6�n�gW$�&=�f�&����O 4C8�q��[��9��`�a*��E��Ig&fpR/�TA�0��Q!��|GV��bڵ�A4T�zPk�`Q��轃|�� �7V=��.y��X�0�3,����{VVVj����i���N���5D���%��̸�qd$v߫/���o�ƭ�/�_�|����M��V%nL�Wrw������o�Z��'�G�#��j_|�|[6�v��4�_�t�<�$��2�\閟��c�K�[�i\����xu@$tu�̎4y|�I�q�@��#�L�3��B��1-�x��B��-������hE�jӼ��nɎ�.D��2�t��B���J�t��� C�ވs9K!�%D��j�t=Cڦ���T.�iV�'���n�vX�b��
Ѽ���p\+����O����hD��]�/�l�|��ؓ�y���D.k`CC�_xX��
F��ݲeބ����
!Sn������J�g9C$:RRR���69!�խz�Ǐ!+��v�#Tۃ��~�P~ۘ���X�r�.��m���ZW*��bcc�i]�5�w��'2��{a��`Ժ�i��������^q?�i'}�{���Cgc	�GD�� �~r��������%6��<�E4e�'ͯ�X^�83_uR;!Өtǲ��n}o�G��΂Ϻߪ��Ʃ�I�Q�tuu�"ˊM����h���w��}O��݉
�/��g'c�S�;��:r���$�\o3��i���IӃkb
�q]�[�銬?��}�T?-;�z��;M�����FFd�QO}�e��Ev�nH��w�wҁo�~~������ȵ�00�n53�9������j���������0�����b���K~�?�#=�?s�|?�)�aL1�aO��,�|g�MN�k�]dW�Rc u���[4��WH�Y+�J�[��TL��;X��쫭5���{a�Wm�։�Ýu�o(&dJV:�]�
{@����R�A�����R�Kd�Y�O����7�Jb ��J�96W����r�%�Ҙ�wyя~p��MU|B�\���Ѥ5���;K��",)^��}�� 7|f���<ް��a;XD��U�{���UdOJ3��.��^`�i����0TY'A1��.׆��U��+��6 �y����>�5��?1��Z=�0�}x�s�r]�������H]�R�6��Yp19O΃��$>�*��g!���PU	�ת�j|T�"f��&�|��Љ8]+��Z5�'��3�z�v����xH�2#�5�O���CL[D�E���~d}�XmLP��*}DJJ|k(����՜���?�	�j{:�t�֠���A�%j��W��ww?��h�������~�y�3��͛��M��K�ن]v��c%��'����\U}�����`�M7D�]��f"�˼�݇��d5�8�`�%[��i�ʞ����G�r�J �����d��,X<W�ݓ�:�X�(Y=�6r�˧.�'1?q8�Xy�*��>����i�Vw�]o��H��Z?;�S=�KMn%6��-R�>|��#�����1�h��w������n��YY p����0����S��d�b(��~$����ض'���iK�E}[Ԭ��aG]��p��s����;�d9 S�F�h ��l!2��5�&wO� ���yc��y��#W���,V���@N�R��(���5�/X5I�}��uk\�n��S�a��Υ�I$��pw�O�E3�ZY"�us�Ɏ]��*���Y����,���!�m Db���^�ٓSe׮�70cZ���3�Y��j��HϚ�`)p �3td	j���:BԚa�z�_10�q������I����[^���}�(lhG��dpz������ �T Xp׾9$t�Q^�%|BE��	��vC$|�BB��\�\.���4���G�KS���D	:uE��_8ܳR�z�ﾗha�����ܟ��_�����F\m�m�^�~{\N�Y&5n�������x����d��技�����'}���Y]����=A�7�?~��p/�p<����ي� �XT���b5�����Q��U"o?��W��=6v�}3�'"���u��vҎ:�^,���e�#3��6�@�_�4Ϥ��#���v��	��D�!^��ߏ�#�2s(������^�l���6���E�`��Z�F���~bApҊJ���B�:���0˭<\����
+�	S��f__2�L�G��Եi8B�~<��j(�a��ۍ���
t	�A�t������Ql�?���;��T�(�~����ϟ�E<77�:�]=׫�Ϳ#"�;㳳ď6�O[���ٹE����$�Aa�s"ͥw��4S�������K�Au�l�>�w�r�^ˈ�n�a�
W�&ϡ�qv���h�%��C o���T�ͽ�#S��7}U�w���%��9Lk{NE@�IH�J�s������v`S沊��V��mu�[��[Ws�'�'q��b����lVū��'3Rd�|�v�oو�9�sʊS�Sbr}��փ� �./	ˍ}��w���$��@����+�[�`�����0wR�U����u/� �9ߊ�����]{rp$T
�=��?���<w���(�W����ll�@O�bу����V�6j�
	���P��uW�r�������j��ٛi����:�5���v03e<I��雿����9�:����r�TJ�O"p�k[����X�MN�}�V��>�T9�a��`�|g�e3g��%�=J(��������n-�&=��1���Y�:3ik;�XX�'��ɿTr��u�;��ם�3���ؤn�JG�ո���������k��.k=�-�M
m�%�m����<'ƶI������!�����z��w]��hڷ��m*���h��Ρ����w<!�~�e:}��UL}5|_�Q~�1M�.�f�-z��N�c�-�HZ�X(�m�u�lq�����o�W�%�_h�O�}� 	���܅5!x��">`�쥋G�օ�5X4{8B�jɾ^�����.��Y�G��KO����̝��4����:3 ���Z�t�M�B|"��t��~�v]�Q'�Z����mb�9��+����)��Ĩ����O<`��ї��ېQ������`�HT�7��1����V�J�Isr�7߀��׍NA=l�58�ۖ�E�k�\J�M����i� �c�%Yדf	���$~��-�K���^a�f����i���}��faJ��?<R2��x"��T�ڞ�G{5�ܨ���hf�r�W\p�iK7� �*��`���y�������6�F����u��'��;� k��Y��D��QP�F��mZ�K�LReW�0��iaϽO��)�9���ā�Z�����>a�Z81�v�=���x�6�! �ɲ�`F�rRE��IN%��7�SI_qUٞ���W���2��1�5���ju���+* :���-��g!�q���.A��A���f6I[����<ͯ��U�ְ���_-����z]��s=̬Ad7՟��,�J�����\ �W`��ҷ,�.��bO����v=�Ή!��fg����v1V�a��<���E ���k]T7>혧m�����L|�e+�%��	��	���6��2b������< 54���a!H�ǡ���q�l[i��-�zD[�ٝ�eEF�K�NE�ms����8[�VO �ec	����T���\��ġ�tn_e}���g|�G����$��ɫ`"����(�Vi��TD��)��x�i<O2��w�}�QŹ�9��h� x~m8;M��{�Իi�0�W�x��=���sY�p-����!V�9S-�\��d=��WKڱ�7Fbկ����ڛV�~;Y�q��|�T��o{���*����7��W�\��iU�x}svdS�������m9��𨩼��	^%������y趻�
���*R�&h<!��z��i4���.�qݖ�X��i�����
��	B��� s��*-�,�0C�	-GJ��Igj�AC�O_<I��r�칺�i�/T1}���ȱ-�MX>W�~7���	���4+�B== (�`Y��������i~��a�6�ϟ�;��4~��v������MO21�������ȠJ�g�n��c��7�藏��X����hbgN��l�$;�����7�f@���c7�lI�_{��&Z�}�dp���M�gm�I���s��x���;>f�f��ʏ�3�p�>�zqn����^N��h��B����ل����܄-+Q� �^���9b�
1s�np!e�6�|&mϚCQ� HK�V���H�-�=v�ǯ��2՞=��әݟpjmo�Ƈ�����p�/j��&gf���C����-R�ƴI��;���砱��VX<R0�v����sFh+�OzÖI%ļ�v��l����L#�?M	�
�6������w#���S������]���^�f���\�"HJ��/�0)3��J���dEQmX���GD�KO<*�up/�#���<�`W���AL�������N�"�NA����Bk�O�,�YO������E��J�~��ȿ̰A�\�G�YR�v�U|�E�5��@ n_��9Qבff�k�8����{z��q���{��5w4,�R���ܟ�J���6т�M�����^E���
� 5$��|��Ϟ"gw�4�Z�pn��-�;B
�-I);���&�d���-3�d��j�kof��S,u��b/F��i�0�H�����V��,�������]]��������<>����)u�^Z�K�f��b�F�����s.��7���/���5�6�����>O�c,�MQ��쳼S�9�Bd"9M+����C"��X8zR�",�:�$UK*�as3g�ʰ]��D�s�,9&�	��8��2�v�����I��CN�]D���>��P�7�)��r�\"��ֵkX��Nsj�U�6�Y�pk5S����－�	�<�&��2�dl��qWߙB�Ak����$/�Гc]�:���Y��5M`�	�2�*e��y�X�:㬝y��d�r��Xi$�e�T�@���_���+E�#��p�S�B
a�<�&��vpM�h�8�!�^*j��M��r���`��*NV3N��̲<�oayX����*�>E`Fې�#���`��Y&��3<߂M<�H�)h��x�<���'�j�����Pe!����n�my*"�b�CpB��'���$(�M�E�����0��"�ݣT)�&���n��T~�1KȽ�����93�Imma��p�c�&�+�!�"i "���=n��|�%�2\!rI��n�\X�aaG�8Y+����CĊH3QRS�(���96b�p��K{��j��U���Zh'�Z6F����qR	6q�<u�2�.v3��2�3�����#�b��8�°i�.�i�5P�Ip��ǛD�X�]|��v��(�B@ɫ�F���4�P z��j�7��L<&�F�Tf�J�9�T[3HZ5�7�"�-�!���t����T�P�b4�xju|܇���4�e��(��e~�!�X=�����~ON��I7f1H��"Ե6��y*����^���h��/�{�qRX=�i�x+=&�p�!�.+'y��&	���\f�/��`
�a}��� \�rח���E�����*���r����(�Q��l��"b�+J	��9_U�o#J+T݊�E��744��ʂ�?��qNyn�D�t�^�a)���
��庸��c�utthdY;>�MW遥B��ٮ�����g� ���Qu�5�*��k�ŋ�q�fl���Ί�齜�S������������g�G��'}U$T�v��]�F���h�����D�^���G\��T\�Ȼjg�I�ѭ^�CW`-�Ǐߎ�[)�M�0�;�q�SEp�3�����tX9M�w\�=4���2K�>����l;����T�J=gx�[��k�����_���)Ƭ6��pC7�6=��_d��*K��ʍ�E�9�Toc����o�o��u�N������������¼Ԫ��FIR{>��V���=�f�6�;j
w���`��Yҁ�Q�o�7f�0�F-Ɯ��Z:�<B�N�3�wkf�i#M��uw4;�NOF
	�:��(�(119e�z7�T���『s֓e�3[�TK�f����C�o~
Ж���޲(M�a@� �k:�ӟ�m���a0��۝�����sѿ�4���YY]�W^/�Mk}�����-��������ޏܛ�nW��ݹZ^3yr��GaA~����F �����>�W����Z��z�TO�3H�,��*�Q7��h�ŲVd3	$��Z��ӊL�I��>$x����r���Fy7\h;��z	ug�/rl7���5��]GiC��`U�W�x�m������c�=b~>^&`5؀;\�ɢ��W7ea.�Y�	����]�#���[�����9HZ$
�(%������ADVk___�T�u-�w.�0�j�w�,�Y�����/6V�lŗS��k�β�f~��d�$p��d������č� ��B�@_O�,��Z W}�\QQQWe�ţ�sk����ѨՈ�.�*��It���H<s��1Լs�3m`�\�ߴף�퍳u�[�t�-3T�"M-�cֻ�[N	�W�i�ik%~]=t�;�S�^��V�($����D'�E4ow�!L.�Pwõ�@�W�pn9�)s'�b#{U�IH����F��g�宂Ƞ:�24i�bF���z��O�َ����#Z{��Q�<���ȗq,C[����N����+#��"�Q�r�(��s�R�D���Od��a<���ݼ�����򽳙������1wc���8ˣ�����'��'׷&�p�닖p�(��֗2W�@�Rix�5]w�"�
l�/X��^n�[�O�ʭ^KL���������'`Re��CL�>�  95����ǀ�S��OB�$��4Ұ{�Q�<M�O�}��@��6������Om}}sGJ�k�&i�̃>_ U/�"���:���{S�S�'f���1eW��"�AuG��q�3�uA�'��}��<��,i�~�N펀mm���oOl?��`G�ҧ�I�Vj���ǽ�X�ˑ��l-Pr9ew�Vz�cs�45���5��1��L�[6�VeL�{4��v��Ę
�><�:T�D��	�Rqp��ɚ��2c�EpU�ƉJ�t�%"X��ޓf	�iWyt6�ùV6ǖW��7�ʑ�ѡ5�`�� `t����ۡǂ����m�K�x�F?��2'O���������]{��������S�>wiO��#�$�,GZ�rk�3�
.Ȣ��Ip�H��8�z�V܅x�8��P�&8���8`OޗC�6,�w)�
��k�w����M�����x;�O�a^F�j5gkcURF&��J+���c[���9�G�]�KJb݈oYtZ��/]�oұ�x�N���f`F:��C�C,r��G`sI�0E�4���>���6&$�Ez��ua�ǵwůîE�\��v�-��f.gs|�u���ͦ��)y&\ Z[D������P�}�*��������	�eIGϑ-��z��׺�	���%K�Z�>�\��2L*%��Xuw��+�BS�F�.du=#J���ȏ�����Iͤ�FM~�0g��p��?�"�]#�S:Җ��x�A�lQ����<�"�|�TW��]$p:�0+I1�S��1t�N!�C��t:�V��ká�}T��*K(�@J�(C�PC?��O�Wq�^����ժ�T��u��b����-g��7�fո]-�α�����Z��ߵ���Dj��i�o��7 � ��3NjffFa�_\= ��̛���{�t �|��#}g`��]y�����&��:Ln�1��0����J�����`R�^�1�#���ZaD,��K�dC�<cU�$:��s��t�b ����ge0R`v�>��]�!�ָ��B�g���ZuǍ;��E9k��0�����[��w|�o��o��G;�������*�/�����a�~�'�ϨEc���"f0�a�x_��Nd�z������ң׾�/��3 ��������^����&�H�m�GDv@�e9��[� �j`e�⁙�gg�P�=S 	]<������:�*ץ�|2B���@��5�����ͽ<�v���#F?�O ��1����G��S�=�m��'-u�ԭ �J�������jm�-�۽u��E?v���㧥���i�6͕����-()����Q!`��͟�(L%:�R!_���\#�WmnT�����+k'�r���,#"#�O:�ۍ�����Cuuj���jޞd&�kh(��5YvMX�|죅�� ���݇��Eͼ~�e�N�W��#�@�w��E�4Kl����ov%44t�&*m�u[B�Mu��L�@��dN4{��L�@��eFJ ��o�G����k���M�n�|}��rI����2�i�!���2Y���2e��5�T�GJ1�R�"X�߽F��u��笵�`��d�FJ��X�	*�z1T�U��EW�S؄����?t�l��f�D�v���
E�,�a�ag(p���H�x�܏��.�J�� +��j���M����;���Or�����篍��8�jS{�Z���$����T>��u�6\��k؄`{|�\�������b�}�>�`/_N��2T�j���%`��}��f����¾����!��؅��KU��8����2�:��O̥�*����ED�2!b��f֜��M�[�~�x��L����� q	����0���O]⤳��~׿;�_���wJ�\N�W���a=>e��P�eh�o�F���^/�� L��oH4P��$
�eU)!\�M%Ŕe)� �8�rt�k�?W�\Um臔���G0��ue�P�l��ٵ��Ժz��'���S�O���`񓶁��P��h�j8�����x{�-�B��i��Ձ����X׏�(S*�a���I	�E[���ź���4@�� �<Jħ<���d��|�5aD7q��Z��9����Ш{�������v3;�{��]	S�l.����?�i �r}�����|�\���m}��M�0kјwAu���s����\����V�{*��u��	N� ��6�:e).��x�sh^�Bh�s臬'�&Skp�1`o��]=y?t����y��ڻ���\��R����ܠ$�-���Y4u3^}9����U�.kL�=M`�7�ӨŃ�p}mm������Ղƾ��\\̠}����y�}��!L`�~m0�fqǕ�+H��D�-� ā~8g;�d��O���4RI�p�+q	�k��G���5nr��T�jf������:q�0SKtB��T�e�3V�>�jc<D�y���	e���{��+��B8�|�i���0V���� �u>a�v3<rU�x�R�K�h��l]�~}l#�	��+uR�+�mK������T����\��
�ٯˑ]���"�j�l�6�D����nj=i-��r1�S�G�W��fx$<���������.��33\�����
�g^Uo<P)m
�C����^I��8��N�x�����"3��
���������<�Tm�� 뜝6��A%4����
�a�2�c���+���sD�^������}�����\���q�ҷ��;���:�����U�d�N)���9������*A�O9�?g!�$z��}�/����?<6'A9�)B����:��ܼgI��9=�r��OCv$����r#;t�4(���}g,��)4I�`�"K�� L�sw"4�4y\��ql�s���?�c� ƽ�6x��D]vs�;s�n@��y���H�Htk�@/`�pW�k��UM���8��e�ԛk5��:S�z���]o�^��fO����dt�Y��=`�p�+,u���鎵�����Jh�o�p���W*auu�����5���S���`�=�ύ�Y�?����P��~5q���L#4�ҲuH��#̣�o��5��Zvf7w�EG4m/�hq�U!#��.�p&k$�è<u�ģB�6����\�ث��s�'��=w�����I��Ƙ|���ר��dY=n��d
����c�0.yM�N �r4��0��+�iM(�}�^���/�S�Ǔ�]�>3!��_�R����2��G�mʩp7s@���%�m	��Ǐ�*���^ [s뾖�	�����76��O�֌�p��G��ᆿy��{�h�~��ĭ��SUyٯ5y����P#��Ȉ�l�zD�nKCEiM#?䙊�S��.y��>��䲽I�+'��D[�\0���B��re�N�&4wT#�U��aʝwonNO���C�ﯜ%�#]������`�FR��":�XZB�4$��B^Flot?���u��x~p��}�1��oQ�b4\w�@C?	��aO�j�>��@u���]j�9g7�Rn�/�<q���KF{1K�XZ���g� �h����q��Y=ȗ�#�-�K(�<8�Y	�G����o���'�p�r��|�-T�j�����"u�'���C=k �`����(8s�$��uuE@m�s��%���ijn�Dfx;�K? z�zͰ�RH@��}u5�̹sG<�d���'��;�6~%\ztb���  S�([�Y޲��f�wn��|�Z�f.��R�� yQb��LJ��<�f��ZA! �r� m��/H�	a�e���{2�~Mg$$]Ꜣ'��Pb��P]i{�g�N��qP�K� ^�ۯ�Ox	nQ�
�������#����y�{%=��������<}`D���*�j�J�]��wf��؇��,�7/�Moe�MX��,V�ط� ���(�a(xӲ,�y0�����k+���t{�J���Li��2`��I� ��	�ښ?G�g�(U��w@;EjS���Z�<�|wJm�?#W�b��{�''m��`w)[ȳ����c��#!�jI�X�ͧ��ҁB ���y8/����N_Ҵ4�!�I	,�?�z-�M$��gp�W�V��'�}�0IBdN��ޔn����DNf5z����0C5`ڤD�2�Ż�ʧϽ��W�9}a!�tdE�s�k։a_N�@�b����9��<'!�v���Vb��Q6%˾���x�<����)�o�u��:�tE�z��k[(?	�c���I��VNĉT9��[���9f��!9�G�Z��n��^� f���9`��l����n��������V�%�W<�¹t_`> �o������'��qRe�4��p�-Dv�s�{Xuସ~��s
.��^��J��+u�VuV�_W�'���'�5r�j|FҺ>�_O��`>;S��+�4/.F��`Ѭ����e	\����\�^�:�4~���/������. ".��1D⊇K)ѩY6o}v��1�T���\��%%Ά�d���;��K��2�v�4�Փr["�i����z��W�\����l ���$�pf"`�GY�R�1恫�[���>?���9��TqeY�'#�͈z����ԉu��W C$� �s��G0���!g��V������W��:g�W��Tr��(��l{���t�H���i�Xﳿ�O�	Db�� )	��m�B����g��#~�Ԗ�1�&^��q�9���I׺���+�G3���-'����:�_�nN�-�V������1���!s��H�OdL�<� ���(W��ts��`���t��x8m����6��Ʌ��J�i�>k8;U:����^w���K�o�pj֑�޵����<���-���GSf�y�8��$��������1��d��.)h�)��y�Wjw#^�zՂ���'��K���c@U1ft��#\�\�K�i7��:;;�R�9E��>��i��n�A�4��r��bI�>@V	w� J��Y+�2b�Ļ�/��F
{��jͩ�&��6'�P�Y��n��e6H�\�x�����n�\����~��Zk�p��2����P��D<�շ�`���F�=��
�a�^�m���4��Xd�5�w�1Y��{�O�cO�W����Npq��j5�E=�S ���R^�F��6 D^��{��#b\]����]��U�/�G,|k�V����q���iAn4	󝁱����ʐ�%���K.p�w%c��J�0�����H�'$ �v��O�v�Y.�j:Y��?q8�2*Y��f�_*Y�-l�J�cV�w~���r�mk��`@k��7�ˎc�	���ؼh����.˳����1�p���
���H�AI��D�1!-
��Z��O��;�M��b�/\�Z5�t�����5d�-�KŲ�
!,����4�G%27�U�c[D�	NT�X�	ɝ��������X���5T�9�>m0yN�8Ժ�e�'�=���1©��B�w��$?e��P����Puu^U�(�H�?Q�'�O�O���(1Q�JZ>�I�;�P!���Y��,��̞�������׉��vQ�����Zm�Q}����iհ^��
�7��`�9��tx��NV�%��R'���T���
��,�R>竵LN�i~�H��lR\���t�[����vb�[o��0hr;�_*�	�|�*����*_��B�_8E���F8�$��a�){gk1;ƫ��"�}g!Mګg��;w��!%b�Ef����:�$�������8�U
n/�hXo�������8ͽ2�H@�VVW�`�*�^2B$�,Gj���l	��a����^֛��;Q�o�D� #��Tk�@g��si+Af�N�O���G��dzp�_��늄U�bT��߽!��A�'Ud�N(}�"6��%�%���R<��Q/Q��\���٘��ۭ^^X�p�wo� ��wL�~ 4K"�+ǃn�i-u}�����Ez��e��_%�%�s��
��:�=����_���w~��"eF��+�Ӯ�z^���W�����b!Wt��;b�,� +�w��ׂ��y�#Ҍf��&��� ����xt�G�()r�$��l���\��i`�D5��z@��w�gO%�vE�'&U-2�pN��vTF�Rɸ�+|0�C�Us�k��/���6)�'	'f�c�C��;^3yv~O���kA�o�
~&�r�ͮ3��[���ٻ�t��P;LtO�,�����{���p���qh�:H�+���i��9�9��v.��w�="�,���KPv�O�iZ�k(����]�z�^[����DVu,G�WV^�˿�ELo}Jgl�(o��R(f��~<`�Ԇ?�*�8�-G����w�>�/N��d0I�=ԍ�?Ƹ��g�R�9�m&� @B�%��d�s��)q�#_	VL�����TsvU�I����U��9O]Jdd��?ؖ������G���X��κ���bd��-��g6-�k �+���W:^�����Dx�4���U��k.F{R�ǂ���o˕7sN[�(�����������x�O���C��Y�Z��]_0ؙ*'<����x5����.��}D���Ȋ,7
"8 h73]��S�4�'e���|������B��~�\e"t���N��UŮEF��$&Z@z�·YN���cU�'���k��0�;�b�u�Ⱥ;\# �Uc�hj���/������4�ۗ
�f�N�<�U�,o�6yThU�bu���Ⱥ��Y�q,1��^�Y���4*�eo����I��?��i��8�������A���>l�H�[�˔DGm�;m�	)�>�Ymf��}3��F��~Q�߅L	�����
H3q���M����v��Y�~�ԃ���h�f�3��#��U>��H��z��w�եjXWq�8�Г���`�R�{��F`���6!�����_<���t_��]tI��A�d-&C�:ˑLHi��y{(���5$g���M>�0E>��f�����,K����f{|c$3��
̆��C��ٯ�T0vӿ�N
��D�zpKj�N�!ჱ
�xdm~{!�@�-4�c��o D�����y����j�*�`�		3�-d���J��
��>m,gϣy����jc2��q�
�ATB���F�k�/�J������#At��6��Iʻ8v6��<%1����sR��ATzЖOgC�Qe%�g��}�ޞl<ԟ���$V*���m�9E��|�Afшx���sv����4�F����y�8�K���B�n!�-! ����롅ٞX��85�*~�����[J�(�ߡ��������_U>�~�ֶ��S�����즋B�aM�j����eH�E~�G���s�Ӂ�.hᏊV�g(�R�4�̚�L����a���'�ș�0,ib��8��j��L�p�� ��P��Y� ��5�M�svNIz����s4���1&���6�Wrk��Q��u:ܥſ0yV�_��[�v�f�����U����29���eCť��a0Z��7Fn��l�ѵ�k�1{��� l�~/�+%@�Z�>0R��+���G���ꀁR�|>����Y��Pmio�e�	f�
�͛+�揾W0��ͤJ	�Cs<mG�|�.�XTʾڑ�"t��~Yg����=:�+�v�Z�}f>VJ䗢?���/�|�t:���H=����&�8RS�V\�U�<~�|H�d�S�����_l�b��Y���9��'�����0u�Pu�'��D�R!���d��"�W�i�,���nJ�%�(�i,[��6d�ƒ4��6�GR�s=�������l��9�����:�Ϲ� [�N�GЬr�h-�;�����
#gB�)t�{��BY�Y���e$��،�	c'~-Z��)��S�����w.��x@!�o1"{K��G�m8�B��g��R���b�)|����GU�dI��-��>_���[ɸ.�b;�G�Mْ���2Ic=r�dť���zd6�j��*?��H ��m�D^�2�_<�)�<���d������x��2I@)��~��?]n7���Kc-�ݦ95L�� }��]�WF�����&BO�*�8���VVƸ��Eu�GV�b�����:'{(	ۍ^86R����W���{��Qv���k46-uf=ܨ�y��8ӡ9H:���eڿڵy�z��$�!����y��@��D6t	���ESjW�;���&'שּׁ���U���}�������ǭ��g}��!׷qQa��y��Q�����������Q{rҬ3H�����9]epÍ/�ԍ΁&+FG���ߍ��+R���k�5&j�b ݅3|~ɒ&;v�9Bn	c�#|�Q���3�⾎�u�e&�����'2(��)4u�wU���_��� A������w���c��̅�Lc�G�λ߳�8s���\�쯌������rV�B�PJ��ϟW���o�6��X^�ʾ�:���q.�~%(�J�GFF1�a�7�e�-�A��	��7.�v'��̦�c��� �y�w_�d*�K��-��P&�0�O�Bb�'1�|�M�"#��{���!Z�c��l��}r�ʐ�k^m���+��
GE~�s+'^�:R�9�����OY�F������zq���:�*�Z��W};�x����xܕ��צ�k�iO��fU����.1�	Ү��+�z�iL�ܚ9�B��9g�4f~ ��e�w��'w������������B�������9DIT���J�E���)������Q��;�)�Nk�Ĥ�Z>�y y=CI��p�ޯ�py�I�lRS�C�T;�W��^K�ձ�j����ih�ÝJB����CU�f�N�,�]
l�n�DR�2i|�7*����)�i*@4���AoOb�s���u�G4:F�ħ�n�U���Q������r��4w{���c�";�qʠ��{&���z�Ev��"_S����5%"�V�����RY�s�$S���)���2�=K����Guv�JJ,����7E�����t֊�sj������3�S�k��9��F��y/NI�K�������� (�Zg�s95H�XG�˰煈�b2�a�<bp}�5��u������%�9�mz�4P�%���4� ����KN�M��br��xZ;������;,�T���qB��%1��Hw���	oE�:��'�i��ΰ��O&OO^L����F���V�ĩ���.��yk'˖#.\�����lJI�\���h  rYv��N6��fw'u��������@�^����R�a1_���1�'���=�������4F_^��n��������&��r��WJn���i�Ѯ����e�;㌻YB���ˬ�XSx�T��O�=��J�ӳ��u��Kn	�3���\�̓� *��R���u��q'dE�:Ԯdȃ���}u�qȣYKZ�ȃ#~գur��"�2�.�c'�.�z�x���y��*�!F!���ڽo��^,�`��j�9q�&o=�lI���e������kR��%���)�* H�qW�pxD���'Y;R�'R0��!�.� Hj��1[!�5Ќ�G��샻��rf�d�_���2����3N.#��y'<������W\�XA�:��K�-��bY�%�cX�HF<G��֟F�jX���_U��T|�}}�;��6摏ww���&v[˱�$�6�C"O!<K^�[,��:ܛj��5�pZ	���7�|�]H-S/��Y�r]c���S8��Q�hz;�%�P͠_���;��:X/�dԩO\��_Ə`}RKV|��
�H3Z�Sg���DJ�`wIO͋�s��, �+X�w:j^���2�Ǣhl���!�c�I�
L�֐V��>��Sןx�X �t�4m�ⱡs1>6�LC��y���D�?П�)�����JcR���-Q'Ǒ�7�����EE�����fy����7G����W\B�E�Y�,��@��N~o
g}Ib��Y���xeͭ}�|lN���ӑdR�1�j���3w��-m8�:���y��;ʟڭ��黯�K1wL�r�CsPq_�jU6�j\���p 6�9:�9�ů���܇��� H���s@#�cd2�L�x�8r4�xc���]�qu��s;J��SkK�J}�P�!W=�S
� ��W}��I:����c��<�7�5�o�e�d�&�i˷=�����ƛKg�\���o� c�ϯ\���fy����5�Z[�8�+�E���1�]�W}�0�/��	x����h�72O|d�S˛���>�3���ۺĆ�c��Z�<jt��7����a](��Xݜ!ɀ�hA��i��1cy�.�#&&��B3%Z�4	G���r�z��EC ����49%ǒ�~�M�'=�����*V�����F�� s�p>|#�Q��^p��Yg�~������}K{����Sa�Bj�Yݗ�b���RO���{7Q=}���)Aɳ:�Q6[�|���'5��o��i��� ����7Аw���wR�_�����}TK,&q^S�!Ü��9pES�%M�< 'PS�����>��/�v��0�YǷ�},���QG^��cRD��n�T�(�g�( =#AX�Q��|��U��Z�|�
��]}'݄ލ��x���M�:��io5P�𹲗�g��d��� w0��M� G��U3��ǥ���){��ñd�s(�zʹ'^ ��BO��0�X,D���i5���绶��GA�P��m+�u�m���N�`u�9��]�t!�]�L)G�_0]Q!_}��1tW�)H8l�jʣ�d���L��P���H܉��'���=/ZC�~�i���1�?<�,&�V�[��'��Q������=�j��,�:�"U�/��޳�5J1��� 	~U��;�2����Ȇt�H����;s��D�_޵J��B��@R{�Q�d�y�) 3���I,���< p����nk�Gjʔ(��M�O�$�*�cȐ!��H�`�%�T-��D��y(S��sS�K�hV	��%��ЋA�־�-���U{�?��*n�簩I!���[�ISj�/2�umrk��L��<6��︨ޭM��w�ٗ��ř��V��B[��a���dJX���/c�\��ȩ}1�=���d��[S裓y�©��'yIƕ<{����I������`My:��*tAK�2�$�U�(�[��@�O�i
�uN|�-a&.^w�;uZ�Ur����T�0�6�pI�vU2:\:%�����dڶ���v�t2R�q@��y���{@���lиXL/kG>:+�Ur�>(t�-+����1Ш��KT'u]�nO�!_b�;�*d�B  /7'��LJ���ʚ^�=�ah�r2��8�7�졲�;� BD8��HT�I���u ��e@��H��+�u�2��9��`��Z��Ȗ�e�҆�wS�a'�dƢ޿� �Z^�θ�iӵ��v����mQ�Y{��%Q2.j�|#��	��.�Qz�W����41�:#H�9�S�E|������ڰS�U+��1��)(T�%K
�Y��Hc1�-Uf�@=Fq��&R,��_vwk�"���H���j�����GF�_�#���v�������dN���y�h��v8��_U3ڿ�/rn��z6���
�8�!U_Ѧ*G�7��df	�\^�4�%*?�X�[�Mv<Q��xE����r'o\�ԥa����q�b�K54��U�.ego9�L�Nc�b�m/�V9_����hHh�=�����~���0?$�bI�3y���aZ�o�%�,n�#i�oڊ��3���9��RI�[m��:hAKO�=�EĎ2���~EN��v�X������x�r��C�F��Ɔ_?��*t~o/Z������wW�x�PeC�a+����m�X�T��OR9�!@�U�W ��&jF �N&~Vm����tH1�"B:��Z�	�Hg-�8�P5�Xkٻ��Y~�;�ˍ�O�(�U,��:{ǋ����!>��g(FE����c�U��wWtZ�wt��ך��O�=����*/ k��͋d��pAJK9{U1 �͔�z�GGd�:�8�'�8׵X3�3]D4��Y�_0��N�����^�����x�ġ#P�]�Y�s�7��	�,���k�#�}�I8���w�'^`[9Zog�^���Y
z��	���rm2�u-'DҀ��OY�J�F\�;E�<u`���h|���`V����b��Vd�$E��5���MB��8.����~/�i�C���v�����L��j���2�$��g)Y,.���Q���Еgr,����k*�?�,���-�4K'itP��F�3���������V@U�lrv�꾠W�� <ƍ{��B����Z���k�b�\ƹ����eu*d#I8���L�Ŧ�c(�����!޴��*�3��ȷմ�_�$��6gY��$�Ϋ�ǝ%��?��I�boB!u��
����ne�`��C_H��R|�m�vm?��!}ڵ�[�c'MqϞG{^Dd�w	�Q(�FҔ���)�=y�m�5��(a<� .�������	HD0ż͐E�W�`s�Fɱ��R}��f��qT�hq.����A�Z��u�wG�<�0��iTv�̫��3��R����Ω� �ǯ:+	3����"|��=�`���`��j'8$�� �Ԓ�A������GR�*oX'ʢc�����e�����>��!� �������aC��|�2 '�(lx}sÿ2�V^����Eؓ����q_���4�V�����T[�|�*6uZAɦ��C�t�.@�Y�L:;�zx�����w� ���V@�v���ax�S�eS�P�K򤰜YjQ>���ePGx�]\򾯲)�W���Iꝺ�a1��<��
8�p ���ä�>ÿV�J2�!��j2�!�)P5FB%��J�:��<�2vo��ku��Y��Pio��i���C�O����>�v�lJ�c^m�� c Һe)�-�"Ů�@ڳ��CG�u4���G߂}���/��ۯi��b��m3]Z	:h풧+��#~��ΦUpc �J�(����M-���L����
�o�[0�2�`���:��(-���+%��#s��eB7.���w�.Ze�޸����ikO�.z�I�toj��/,�>M�r�-U����GrN2{� �������^���*$����f����o/�V>>d
L�i(0;@lH*����,�"J5���cQH4ܝ>d����3*��V+�a���{��4�S3��g���^�?�ݯV3N�fu�Sdc�_5��'�ʰ+8(o�>���3U�5R{����Թ����sk�wl��S����>�X��{�X����!�-�0�� n�6�q�Pٻ��L�"Cf����z��7�����HGs_������`B�d��]f��]��b?�Om>�T��l��ԉ*��[�&�YW� .{蛙������}�e��y����q��V7�f5Zm���Jܛ��|�Ϻ��O3o	��U\��3f�/3��/���
f�/�/����C���/��'vۘ�K�d��Zf<nME�DweZ9̗7S���)B����)��)E�[7�9	��E�P�˄���:�$RI�M,�s���<K�0�����r�F\s�I���C;�_8w	l@� k�J4ָ�>�M^���B��m&�	K����|�ϸa,r�շ'�;���s+]/�%L��d�(c:!� ��?II�nƸ��$�/斒Z����d�� @�ewX3o��ť�a�`]:;M�<�5�<��� �ҽ�i�݋:E3OC���H�"aZ癘K8�����v�ޔjp����E�wc��]�ȵS-c|���dV�Q("���p�s)#	��'��\����%DW�K��|%�ibκ{�U�﫾K�Ctk#�ӄ�4fw<��4QZ�;#����:�zbq%/:�*"	qB\;����-��1e�锓��]+�8e��]m�GMժt����� ZvO�.�qVhM�9��ЅoP=]�L��� ���k���4(��?�n!@�W��!ŗ"�l-�M�}��Er��H{WOM��S�A��F��*b>�t�j�Hq"���I��xP���sSu!�P�qI�18��8u�XPl��$�yM�K�u���w�d'C�J3�2U�Z��X��;����[���ӗ���#��mS�4��`.�WFP) �3���:�3]a��1�C=��X.�!̃��v��7�֯���F�� �6c�d���|�8S��2�x��r��'� ��1ٝ�K%�RU���.�u�i�W��Nۺm�2�f��q�_�sk�y�S~ʀ�����D�l�|A��ޜU���J�R��=K�@���;fW] �1d�(��CZqz�!Gx=�0 nw���1@.�:��a`8|nC�7���n�)�8U�9�Ԑ_���m��#�B��W7mAod3���g��� �d�ӭ��[�~��-�(x>ܨ�p.�3Ic�de��8=p��ҙ �R�t2O��J���>�'ט�zJ���sU��`�4�Ql[C���`J���w�����C_t��e�l�E��+Ů.!'>~DLզ͠�4�z5�� ���x�j&h��
N�h#�m}W���H���6{ g
��G�������3- �ؘ�6�/������I# �D^��z-q7J�vC��(��|ۼ|6����'=�}'Ȟٵ�����@�#��;��J��N�Ψ�Q=/z<�����O��/�!} �J�P셠s�v|�W�Kڅm͟~Ff��Ev
��C�n��#��ۭ�/�Z���¤�'Zc�o�����`����
����^:Zq����^br_z%u�WQ:�l�s)�f'eJ�9VI�ӵ���S����q�K������?�*Q����Im�����k��p��w7j*B�ұ�(���!~�G��v*���r�"�����������5�m���j��3��-ô�@��p����a�y�+ɜA�K�������	]:��̮&�rÜ�*�� ���G��&��� �9��e��6�R��L臏o�8.Q�R�M��"L|�]�J���y��G�5}%��>Ⓞ�g��z!��Y�e[ ���yM��ݯ31�g�<��mL/#(�W������Lq�j���3�5z�i� ���^KzǍ��!�MC�I|C�R�Đc�1��9����ڌY���tPS�'��B�C���k .���76�+:�]	z遤����� �LO�$*�-�|��n�i����
�7:+��{��K;�2����SX��Z=+84���nne��,�bl���ş�C�\]u&�tZ����>�݆�?�-ϋ�g�e��ͫ<���d<��:����/|����
��v��*0";��Pť֮�!D5hM�����* x�Jg�:��9�����F�=�}�Y$�B]�(�k
�o��PI�9y��V����[Ex�/:���3[�cT��|J������$G�;1�����/��@�ƀ>��Jd��K1}�U�.�W ��&��s�Γ`H�x�i9�f;�\�Y8ӕf�<u���l��	*'�)Z%�B�8�ߣ�ݏ.�Tx���5�ǘڜ��,+CY��c,�/Jp�N���r�-��7��VOb�5e�S�[O�Ɨ��~-)����i��)s�P"���&n���s3S �iC�R��զ~����_2�ƐZ��|����d�&n�?�^��X�\��{���Ǚ�k6"�>@ɔ{D��?�I�āp�W�&h��XL}�sJ·��M��"�����An����U��=��Z��!��WU<"�V�ږ��c����x�G��gE��|#
�|!��{����~���뵤�O�yCX�`��̦�}/�Z'���"�$u-�I	�jn@���VL�d���[��q��/0L��h�{�ȁzV��g�n�Kťa¶���t�$��[;=�\�qח��gY=:w��� �J���E�_�V����}��Xl��>���SX}�Q�u�wA���0[��𔏾.��V�ǫ�<-0ܮ�]����=���9!l)��S�N���J�o�[W��朐�aNՍ�vZ�#&�F�xA���,ɱ���]=*뒪ő�J>��: ����Tu|��9q���`��lċ��>�,�~1
)�K�������֎y�)�S�N}�"N1R�rfi#ūzٟp��@���[��[��®��+k�L��;
�0�[a�m��=���1R��� �v:_��2���Hf�Ի������l�[*j�r7#�c� Zֶg���Sf��[�`<���Î����ij+w�/=��l.�"�u�2�_L��M���L�	~�����sx�~ϵ[��ۆ�Q��Q��
�����7y�x/d�nxR}�>��5��ߖ���WѴ׃ԀnIB�������k(g�w���ʝ.��Xۘ��8�en���y���*��#K����wɳ`G^�T�U3��K�I�S��/���6rhor��?1�EJ����KY||���ÜS���G:���f��隝t�$�u(/�֖²��G��r��}Վkn�N����
�Nl����� o�Y[�M����O/�}[k8�6��kq��N'x^>v/�G������ȷ���8&�U��
'KW".�CUi
 ����'˟�,KO�=9h�x������>�w^���ބ|�
�>�w�z63��СHr1Dނ�O���g����5ӾAJ�-�a�`�-Цa��z���������?k�eKQ�&��?�7#��||�Q2����zʗ��l���4�@R|�`}ҕZ��G�񸬄��I��G�.�[��z�O+MI��R͛/a�MA�(f�P�����Z�����3��/�0��جv)r[J�����������B��P�L!v�߬���"|7��`��k����>uU��1E�t�ײ8!�K����~�t�
]��ʩn�X`�)���(t����% ��1���B��?�m|�o�K�i����Y����3	6�\_���5���*�;�v�i)���JzZ�vN��c���t�[C��h�aj;�r�����|�O�� �`��t[6�Jy�<�ZE���$�\=�I���;"r��{�fW���ܣ$Z��O4�j,?���Pz��Qޝ-;�ga���q[�fȾ��.͜k���BX<��}w>��&�2���5?K��7�h����t��]�>D��r? T.�Q��SJy�AY8b����#��S�TDTĹ��_+�@��ѻK��z�Sk���OB�ܭ]� �"c& ���Pv� �Ũ{�	����	ӕ\�
�����r�<�o�{�4�mI�93�,�b�,�� �߸?���Q�5J0d��ÂW�� 8NP���i�؇�۾��,T�F<N-g�����:nB>���-x6v��E/��-`T�d�	��8����*��:���\`�}ʕA��ȡ�r���~=���	K'���XՖ���8�E!Xtw(��5�q�4�����|L� ������Xz��Ɏ�^�-�8=M��N@��^����P`vN����W�� !�	�����l7�,cd"� �$��Wa���=��e�n)�����A��<Qn�vӘ~ӍAu��,i2^¬MF�t�%��B�@���3:���-���f�s���,�F�N�q|��v��M4�|er
hJb9����2ej��lDک�������9k�ጦ0�+�Tg�(�x�͹�<%���WC~J��4m�h<�}�8+�<פy������܉�	&QQd��*!�U�� B_�M�-K��ݹ |~�6��>�����s�5GO�ޫ������#���~ML�<�K�����H����`�+�,�\�絯�����;d5
������{�D,���T����Zr%���z���zG���ϟ��W}�n�0�wr�w���'{6��&g@�fP���_Gd���ܴ^�}��������)�`��l'��Ѹ^������a����!"
�j�Ց�W�vV:Vj��
'�8!.���0�D�T�f�3y?�L��kF�uu�fh�3��W��0`#�pB*<ʶ7Ry�A\^��#eo#8�n����#?_W����v�q�V1'گV����?�|% ue,W�"G
2ٱ������(���]��u�_
I$^���R��W��q�����*��J�mC M>Ɛ8�a���hy�} ����B���_�������Wf��ͮ5|"^M�/��;&W��вh]Z#�
b�Z�^�`�I��eNX	��߾Q���sS��/��v����f��j���a6Rf �HyA� �\1��D�(���"����:f<�`����"i"��^e�	]A��^�0Lq�X����2�RO��t�bk�+
�ys��۪���!��0�����!�%������ʊN�y?�
P�D�����}�IA62��LtV"n^��S�Z�(����(M:k%S�:�z�&}ok~D~0�j���w��.�°V��h/��x=�;q6c�"&<�*����߬k
ɦĞ����_�����i1��`�_'�`�r�tM!��[��3Xe�\��#��PzAD��g�i�ݻ�̌:�,��ЍTm�oTh�-u0Ro{jm�,3hxA�	��4�������#�������\UM�{o��!�K�d�8JR<N��%����ԡfJd��G��#�0��x�L�8����!���d�������Vn���#U���w���p�k,\����hb�=�z���~���S{��U!���O�Bx9V��c�uN�yh��'�)������О:�5D��.w��h;N��8�j�cUsP�7��D������
��߆���a��u�F��ᭇx�l@��e)�O*V;o�Ǚ�.U�K�����j��Ǻ�4�\o�f�)�����>��I&#���)ǒV�r���ә7%�U�����S���j¥P�9�Z���������]Nf��:��[m����FDv�#b�qU�ȉ����g4#$���Q��:���=�i3^�Q�`vow�t�;��E|0�W�13u�< jq*z�ۡ�<�ұ��zHcj}���X0��^�(> ��Ҍԭ�� �I:A����]�c�Yg_��>���x�+�X�	|i�<�M��U9U
/�<]6`��W����R���F�����ڿ}s��	g��,x���IflT(�ǳ*�uP����Y%\;}H���i,��m���v����{[��Q򬥷J��Y$=`������O��K;4�/"��fW���M�>�cj5|��k@7SW9C �3���_�i��l6����<T�F9�q�+q/[3'�hf�gFB��!�U[��RSy���䨡�.YvN���f|_u��8<��a���e��m�<�B�ɟHi���F	���i3�՗�lq|�f�|PN�������7��2����?h^�܃r� �>�{ԶՉ��g�zئ�~��eiO���ɯ��@�YثA��[���HYʤ�}S���o�9�¡;�N˸��s�Sz�|�:C�i���a�x9U}c�ט��p	��]������]��G@ ���-��KKɤ+�nm����E�0���E�:?|	;p��*sԘ$�q�;D;���Mԍ<���͹�*V�D��yvP9�����o0sV]����S����mO��j��\��{���X�p��u�~���5eee'�%s&�8��ಔo;�S��^Ijy�߆!����� �L����ƐZ�� J�G���ќџ/Gφ]0Nn7�N��f\(>���wo��4�����tQ�R���N�\�{�Wӡ(�y�)�Մa��P:��S��'��;��,t�3�U�3�FQ�?`^g�o6���on��1�Ϗ�胇{m���5�74��o��� oV����p˼��T-��>�������&(�Յ���v>_)���=pvE��n7��k�H��]�l�k0i\g4Zo ����b��N��e\��8��N/�g>T�|�y�KI��9�e�Z���_�N<�OSfN�G��ۘ��_�9��KPQ癷�Teԩ����T�V� �S�2�3��;�O��9�>�&1>���{z�֗�M������p���+K4PL1�聭������wQ%y���P��<a�wA]bP'��Ϊ	�ȉ������ڈ�z��������E^��(I4ފ��Π�CA�۠ 	�O�� s5N0�,th�{�)�$��&���*b�#)��G�Œ�ti�'s��x
��JF]��Q,cu/����%	S�cQ��w����a�d6ɢ���� �ր�B3�g�籆�$-��aYڎǪt	��}�mS�N�Ip�a�)ߏ*�ƤN�a?��v�������08U����A��w*�9�j��ob�{���q�	2y�Y���̓�z4@!)���3�s��^c23�Z�f�y-N(��K�R��:����2�%z������$ ��gV��/�,�P� ]ڌ�Z&q�����+���lw��l���t�6������N��a�L���ޞ���S�g��[ݷT#�'6unǍo�C8�<�~�I����$��e
^ƪ���H��SO�Q�HA���������"�����s���!�:m�� }���c&Q��� a�s�@�Q��[���pE,!ɼN@�x�Z8�z��,�U����?m��B|�4���6Qt,�wn���e�1��W��}m&!��������S��^������H;% �.=��40/�ok�vp�m��)���Ee��^p+� �V9�iSBp�@4w
g>�J�*��ix�8?q_��z$������E��;5���W͘o�e:FFn�!$���F��y�^��[� ���yn�j���_��p6�C����L�;pA߁�����_wಾ+��/��ή�S���b���G�G�\�!�_����6( xߡ��FA~Q�I��?��t���X�#2�p���sܫqT��0���#Թ5��/�V���xr������O��z�JG�JB�k��8�Y��Un,(S�����q�>�Q�׷�W_v��҅�Wmv]����p�����~7��n���k���UNH�[kD��=�W[���#�̢�p�@�u��qׅp}��F����^��w��E�hJ9��<�W9Βp��amy=j(r⥥^6�Ҕ�R�^Џ^���6x�Y%k9�vfyx����>���R�(������8b���
 $�;�ı��q�V���
N3�Ő�D��������0�@�*��Z���-�V��!"�)�u�3�̬��<Lb�(����= �����4r�E�������B��[���2-@�6�c�>;��p_�;�����o�:���$[H�k�-<K���
��<��)S�3�^ʀr�8��љaL�f�G �p��-L͜CT���'q�a�k��q������ ���Q@��m$8��$����5�ʔe�F��Y�`�~��q�㭉a���8�K�X�&�2-ӗ����3:�������I���o�Q�P��g��^i�,�1��͍��-����5��51!�A~WM�c�t�pteS�F�&$�5z�=���F=�^�m�U��\ރ�Y6�&���p��b�U�H�����H������er&�����00�w��b2��PX� ���e��yDb�E}ݨ����.�b�7pdW
�fd�\�\�~�7���3�TJ��$j��7:+��$�庞Cu�Q��Ҫ;  ��̐���	m���4��7��Ϟ�1�̈q�{K}+~��wT���=ۈ��U�n!�b���,_1��{Jl��U�~X�Q/'om���M�LmE����~�mL�n��O�洄g]����U�s�X3��	�df�w]���Elt���]�V
J��Hܢ�W��jq��G6���Z�Cj�U��g)�3@"Rݒ�� yڬ����|c;/k톸'�uh���1�p�N'��7jL���������O����tQ_>2@N�NN���*]=�Q���&l7���+O�� �\Ad9�z��� �����@y�@�	-+�g6��I����PR�&���LI!���!�9��)����gއ�E~��H[6R,����籲)��p 庥˚K���fVZ����/�6��&��
��܃C���dn�> ���o�h�s�C���h��5bdddڰm�u��ĳi�,u~���9�M §S��S
�����Rb�j�g�^��L��R�_T�^��/�j��d�$^_��4L+��܂j�'3a$��;�T���эF��i߁�����6w2R˾��c��S�4���u������#��k{:�4�p�5>HKc����s��EG�M�4q8"�qƞêW��o��z"&�]#�o�
c��h����Ġ��P�Wy��_Aj�4���$�p�={�a#�w����w�#���R���W�lK\��U�����d�yM�r"~ZG�t� ��\��m�����_�7�^b=�;,K4��oߩ(����=�NE.J��"}�V�& �����<�[+8�g��?�=[�T��y�� t�ν`p([j򽜐�$��B[-Θ^�>[6��	�v�[[�E��a�T�RJ�<��ob�[�r�M�5�.ne�~���u]���b�i,�V?r��E��n�pM鱙Rc�]'�V�p�k8�����|)�z�ӮT3��zX�z��I�6Ψۀ��L�7O�n����oܸ��?"	I]������-����nϯ������Ks?_˿�ib����i������ϯI�z��#�Oal�j*}K��w)	m���7S��ۚ�>�7;�R��4=�j���*�BŤr�޷<R~���T�Yf��Ɏq����CG����t�R\�Y�	�蘂�~��.���%��(�X�����}�Y���Yb�AЋ�Ft�������C؞���9��bJ��F��f�{6欮��}�7Ͻ����/J��je�c�Fv���S��z����^^%dH��#��n�j����F>�Jh�wH:#z�	 ���"�পc!3B�5�#�0���vp�_#�?�y<d����$S��xR'�������{�7v����s�U#�OB���s�kz��D�r� Zg�C&8��_(�|��Bk��
��j95+DMo,_�� ����h
����JY���]Zp��/\
?2I��h�U@��o�����n(G�����ұ�8��k���TDW�ܝ*aw��Y�Idn%&��җ5%2L�������_S�_�~:.h�^�uM�ה�pXiBR�>;��G�O��2{���k��KFE���5���vDP(���^�]�s�*8}k��F}����	����}#�*��`w�8w�(��7�U�b�3�T?�n@���w^�����{ l��z����!���F�,p�{��qC��0҄>�?H��@����;�X�Q� ������j;�O�:�H��SQ�J��utAmr׉��V�n�P�g�Q3#t>(����a1X�P�p� �`���:N1C���SU�Q,���)EW�8����V���%D9.z�Mk�1�+ں!�!۽�6��$��),����d���9b[���	Z3U><O�R֒�Ch����s��,�7/��������aj
�<h�׆�g������F9w�ޭpy9Ŭu���k�4����-�k�eS�ت=ے����]a�gHmc:j�\�ӎ��$Dr;0;�%��8�ǛYE�-buz2�_mYwkQZ���>�����@v����e����sV�a7
`��Y8�l	��LF��(
�vGoe�T6JR �ŗ�t�<Yq�ƔR�4`3*����-����� �)�S��*^����x�g�T�t�ʭ��l�p��*�m�X�4R�O(pF�;����49n3�ޤZ��qQ�v���}��?�O��E�����#X}y	��CZ���>�4wxY�2��n�r\�Ù}�J�5��ea�w��8��"N>�m�S���/�E�3����Uj'�C��,_�Ip�;-w�����A�}4"T�v��!�-`��y'����oc��-��oV����ʄ9ǫp�z����Ҧ@�d�k�[�K�������J6����[r�,#�&�W~��0����ޏ�J2c�!V����ŭq�`�MI��y�.s,>K$m���%9��k�׉j�a�3N�5��	�[?��@)@������P�ޟ������Ld�p�If����dh�����y���:�x�ؽ�������tZ�m�E$����#5��5����X/ n���}�����e��*��l�nm$��L�B�qR*zK5�/9�DaZ��{��$��W�۞'�˳�r�d�!����~(H�=�&H�X�����&	��^2��V��p����wq�^b'�3��2
��Ug^;�8y6��}]M2N:����5��p|@Mu�Ϻ)�fH9���54��Aڅm>���|���y6�R����pC�0�KunZ�_I��.�p����������|����Eb�#\f��3��ц��I�j�+B�Ƥ@�S���&���!�<��/XĶ�Yg�G{i5N$ܨ�CC��gb����y����T~d�b$�h���?�1?�ɨ�ۇv�!7�}���xAS?̼�*��%�E��n��11��L��o��(���(G���`���e������ m����&�]�Q/�A{))�ŝ�����$VNN���R"�Σ��Bud�%Z�)w���m���N�펿���/���_(C��]���uhf9�B�NS/C{�d�����#�a�6': :q�9xu��%�5G��%l�έ͇�� _A�����(J����4�Q�iA�Y�{���2|���SZD��zb�� u�r=���#Qt�A�@��c_8܅�=�Z�7������c���r��YT�x
�k<�c�sIS!�"��~8�(;S(>_VgKt����|}&hT�MwI���l�$14�-hr�5ϾƘ��xH��ϒiwU����/�&jǝN���.Z8�������1#�*o-\���P�{Tv{����	��8R�Ў�*̶d��	x�S0�'M�>�U� �z�������䮋��K��=Nm͘�K%��L�А�����W�+ޭDa�O���P3~@�Y���7���������)K�-�GaDvBB�lY&e�w�,�}I�(kJ�oI�a&d�ƒe�K����z�>�?~�[��f�3s��y]�<���<������.�zE����uL��J� Np���u���k���s ��J%�ˇ�}}�f�Y䦆&��vI�5�2�Y�Ҷp�d��ᒁBMU�4���>V6r�Z
v�x��6����{���Nt@א������6��T���֩�Ï凗2��qK>^���:e�����Uq�M��t�`�:B�Z�9�a���y�|h���u��q�M^p��8��,T����_�޹T��ݭ@x,�Ā��\��Z\�>�j{���g/E�qO����p��:��ZQ(��$!�x��lmm�(勵L^����yc0���x�K#!v+*��¯ߢ�)u���1k��� w+�@�����N�	�J���u@��E��!�a�SV�Ph��K��Zp����eqp�L���n�\���xP(��>&v���n���:z����������n�_]~�?wY{'_�vZé1�z�
_*��`��k��P�|���P0$|�]��q6�܂¼�k,P�ؒJ�t�� ���[�vv�b�_���,�l�����=��)Of������ݟ�#�g�45�DJ��x���ހn��q�m�?��J��_��z�ޏ+.��8�36��o�ɫ�,�7p��ྎ0��+���!]O��W�b�h$JuzW�L��� ��A��
����S�����7?Ό�|w�.!y�����V%��h�ھ_�	����g���衰y�L(cԌ�<�_[iii��"�R�����U��f,��� ��S�f�EnB�R�ǣ�5��q�0)2Lq�/�n�Ko����k�maK�h+p�,Z6m���hc���=���p�b�O���kT1�c��ePӘfM0���蝆,ߎ�]�P����r�-aE�r�W���a�^��3��u��#����n6wf��
����)�Y��#G z�F�߷:��*���jX��b1i�L�pX������3���C���W��L3IFe�HTi�
�PU���a%���xr��p���yr7�d�=ؕ_PX���� �\
��ү��W��癊LTՍ���wC�P�QH��薹GћhT��7=5����jz`��!x}�؄Yk/�*a�s1Ҹ����
�0��Ƞ�/�-k��~h�D����i ���hKp�J�Rc�IH��$��%���?�?�ap3i�X�H��y4g���:0�v�/  �ۖ�� ��}+Q�e�N2��+��W_h	emb�.-�R+�5�l����k;h#m�2���$��2pa�,��=����/�M��ĺ�v�E7Ub8��A����"��v|FLǂ��`g������c�.di�%`������새?��2���F�������%��p@�4p��PA8��o���j�7|�.�2b���d��lL�v|������#b4���D ��2fb*-Q�*P�V��_�섿ͤ[������mꉵj��5(�t�6U;Q y�sYA��7�pS���@�
�2� ~ �h+	4*��1�؃bI3;�۲�]�n�����R���e勚<��L�)~dz_[؄�}��\��tC��������8�͑n�����ݍ^^��,���� r�J�Vm$�G"���8���/r��i�O�<�<��?@n�w&;�e���C����C��Hw�+�}�����؋(��`�O���4L��WJGU��N��F)��w���/蝆6��C��ӛk=��{�����ɏ��?����9u7����T���ZEJ�w C����ևE�b �V�"�U:o��W��݀����,���e���
=]���G`/Ώ����fY��zq�XM�-��ǿc�d�X��y�]�.�Aſ�2�Fq<��5� Dm������6�=�4Js�O�W�"��C�6�G˴�bi'�}��/�f�d:�eu���e���A/�/VRw<�6ݖ$���Js��q���Ѥ�8��3��,ۈR@���������7W�GD'�=���V��9�#D'�c�n����8��O�[���>G��u2����chx�k�5�87#��U�w�4=x+|�up�V{�0n<�L��Yn���h���0�3���5r2�f��V�=�P	�%���\K�����Kl]�bO^λ����0�����O!�/@{�U7�1����Z�Rp��hcС��y,��wkʂ�"$δ�N����޾o�w�nI�n���/��HA�G~0g��?8�y�t,� �2����T�C�2A�F[;����^�w�w�<C��p�p�<u(�Gz�Z��v�Vn�D�W#��x��6LvTN�@�j�)��H(%.�3ݕš������2�Y9:�v���p(�l?D	i�=Ml�v�#_|�:<�6
�텙x�;Ner�����޻�$-Ճߎw�g���m٩Î�2/tat8K�~-B}1�2Uq�S^^��/c���C}��!��Z���Y3��vqkr�V)r.�f�Ur&����vW�l��a�WSsU��E��
 ���`���e:����Uw�Y
�7�W�Xݟ@�����;�Jf�Ź��9 `�=p��(WVs��7yo�1u���8ZKp)�<���/�'���&TO$EP
X��3+�
�A����ڌ����S��Hh[�T1���9��'�n 	�( @L�j�����Q/T�_Gm��eM��o��(����ɟ/��בR�]��;������ŅE�ޢ��_�c�������)]v�6�~�P�92̌Bc�C=�O*�4�Ԅ�Q���+���{(�N�@ף.x)#�[�|]|g�x�J�Ӽ�ᡬ	+������nq�=�YGg�u�3���_�OP�����P��ip�׽���fj���u��n�eH��!\n�/�c��>*|�Χ���ow�XG+�{�z59ϯ�����#�,N��t�u��:HmF춞£z���X������E͎�߇��n�����mn��=��n½��"���ψKᰋk�`d*�N0���܁�^^��f.�kf�JII�{�F�W??)���X��p��&�{eF����C�a}�1�&b-)�6�"?�3���C�~C�sO�xE���V뻩�U�� ���Ha����I>ژ�%����mvtD�?<2���Zh���;N*]?$³���Po�<��K5������he����������o�����^w��T�>|��H�)ix��{��BB�#���k�{�=*`쨥Df�c`���	+C�zgP���7���R�Z�q,v��r$�&�����/����/�k�b�o�Y5_�m^2���xi���^��4M������ҹA{�d?��eU㘔�=5FށՊ�`^�-C5���Z�L6E�{���0��Rը��W�g�Zҿ��T(�+�<'#��W�IW�h�9Iy�؋S?�RL��<�Wo]>N����if�8�䕤����&��i̔~-�J~8��������y�3/�F29��6�1nDbFԝ�����W�:�Y��ƛ�	��	m���+s�~o�u�T���;Q;�2�C�k��*Aj����P<��+,X��{�/g��������`x��\7��D�'D��vr{	m%�\6��V�q~&ch%@<lݏ���Q'��93 �q8r��8S�;�Y	��.9�=�&�4� �n�íَ�8#��i�U�6aD��'h��ɻÌ����2��v���i��V�L3��:-���s��o�Xyk��+�0���X��ރԃEσ�Z�$��~��]	+�\ݦ�Ro���t�.oI����w)Xzz;��sg�=���})��~�-���c�G,^e���:���(�C�z8�����:(����Au#]���uY�\����B�����J��^��(&����ݿ���Ր�YޜrC���;>�<5�fξ����$�'����vNqcU0ض�m;���:�B����؅�(�����Pr�wt��z3�$s�����[C��r�w��?�~� l�N�51�.�,���ȕi�^4M:�2�Os�*�z��5��C�6O@tPv��)����pu[@}���E�#�U*�̟����ft��� ���$��% �k�ߑ캁������3�{$m��m`�D�HGU�G	4�\�l0�ߟ�i(��gl(�Q���N����3���H���%����}^��yx�#��跾��ކ-  �
�F��Ѿ ӕ���	iy��=%
��8{fe�\C���6�*���EuBq�׫k{�A�`&R�z���ΈC��)fpQ�L��?����7��XU8������{�9����%�LT��#��Jz���Ɛ�^��H����M��f��ϛ��csw�z�4����jjB��Ȋ8�39˘�ճ@�rĎӮM������j��ܪ�(
�"��$9����ݚ�#/E(�i���ق���w0iF��V1� �(�N��i�9���4^��g:A� Vg�5<�(�h�/\��k|EV���=���q�tqk
�G��V��7|����S�0�g}�0�(�x:�5ς�_t|QM*@�/��� x�E?����C�tZ3~#  �?-�-���B	��{Z�)	�v�}C�AoS)d��j�Hě��4�C5�7۫q�DŵB�ɤ�����LeH�6W+���9��'���t�갞{]�L̃j{j�pב�+I��_���Ɠ*�U4j���+�bKj�w���>I�V�Mf��U��dN��ū�Y�}��BB�=,���	�kߨ�*1��tI	�#���P��)�z�֣C�+D}ۇ�>S��G�&�b�W�:���Ԃ�u��7ux�������}$�����k���&�����D�5	/�NH ���_kD(�(�*�8�_�}���ad�X�<7p���o@;mQ�P�ލ�����x�k���(`�Z3�#ֲ�@�ΰ�f蒈v��GH�b۾�l.{�JR�����PE$`�� h������Zq�q8pd��]�Ç����Qh�(��dc�LT���ьYprK��iM�X�}e���� �k=�Q@a�"C��S�˥s�ߎ���ΛpsAL�4����C���t�)qc���t+�7h�Lcm���wX�b��B�5?&4����ku�|zU�%[��${����'�y�l�~�ζ��8�k�S2V5��e]�:&į$]�O��R0���N�Qg2������/P~>(Zn<�}1�I�����v�13�ϋ�]W�9�O����&⹈�� �D�v�1a�Pc�����
�v[F���ZS=j�����jW8H��Y�a�D�0�-T�? ȹo!R�{f7Y�*������as���G]�8�Q@T
��'Ww-R�����fP��9�;����>�~mG*���3�����ï�&�l�T0��b��**�y^���6�ۑ���̒y�O��f���������>œ�t{��zS5�/�HpjKk+ƅ��+o�G���[kR�j��}�Œ& F�����F ��^�4��� m�^�"�4 lد�P)$;�DD���?nk��V���sW�$��	����nа���|�3�h�\d,c\�E�@��������o��}+��=*r�f����_:�Tܟ��<���$�w��)Pc�n,�p3e����?�t�3������i㥩��w�m�@�;g����3�僽ˇO������>�?�Ȭ��}3�rbӓ��D΋�X/
���o�����@�����L�ܬ�L?7��Q�_?��R5kÿ��+����O��D��#����sŢ����\���_�J��+D��'�d��㔜$$��ȸ��=��#�R����z�;ۆE~�������t��;^@3��-//�a�N�`F��_�3{_���םeִx6��$��XG읭sӻ�MdB�)9�Y�Խ��$�kZ%)��d����P����R_�O)zB��*ӏRŭ��w*cEת�ɝ�|5�<G���!�!�tV�(�u{(˷�hd�1Ơy�^��Tæi������3<�N��>V��k���QϠ#mx�O�ܴ?������@�l=N!��j�I>=�FgF=���L9v��4�y��?�m-0�Fi0��!��vz�I�CNݺ/[�F�YHϮ����zw�umk6Ts]�7�_=�X�m�(��Ld{X�h�8����+/�Ww�9M���4���� n��&����8��9�E���"�����Oi�^��
�R��e
c�����}�ddT6�I>���z~�%aBZq�r���SIӋbG�Nzfe�n��b�n �Q�T6��^[�d��L�T\���?Q%1>9�� b��,�]`���Ilå��OD�0!�[��W�ԵE��;���ө|��].0F+^�GjN��r
yw����;K���~ˮ̤�	���y�Y�;�����hqI%�i����d�ZAo�@0Ǹ괄�W[�b�T�?I���xcǵ�X���Z��O�)S+�}[l�rlC�`��������k��b��G`l�#�<�Z�5�mE��d������[UQ3s���'��rPB���[��ӵZ�
b���R9��x��K%.C��~�ἓ+��TyR�ݯYU����f�^\Ѡ�&\9�*�j�9Ib���擇�o�t��.fb�Wҍ4k�i_��m/�~�'��_}�H��c9ؔ�������5N �a���޽{_�R=	S��� p�)�$�J2�/P��G��k6j-���ҝ6��.V��K��QV��A|�*��<�r�M�3���ͱS=t�KR����?f�#���'�]�v���Ic� Orpt��z���9�ǇYC�n6�����7���ӫ��T=����D�w�湄��q�ΥM/�h`/�Ġ;���u��"��[��Ņ�0n*�C�[7��_r��c��U�̪]i�#��b��X����X/��s��oז!�L"�b�8���ݚR��`R��U�w���t����1���� � \����#�?���#t���|��DFl��t���|��� �3ؚ)�c������'�^���r~I���:�Ffi-A?��g;����۱�����е��3��Ӎ,j��X��^�F�#ݣ��^�,tC�2�'~���Z�$'"�k��]D;�z��r��`�z�.��3�!*�Q�R�ҪY��b�Jbq�3}`T��W��Z��"T2.\=Y�����ǉj�{�G�����N6}�y��	ɡ����$�K�|}x܋lr��Z&%&�E
�kٽ/�X�u'V:�Ø���I��j�<s%��^��G�:뚤�6{\|{�QxJ���T�w
t�*��{0���Dr��Ӂ�{��ڞ��6_�19�!��+�5��2cV;1s����/��o������$�(�[#�u95����u���0����x]��8	'�y��� \����U<�O`6O��a�z���ʪVP��B<	����U����Gh��ABڥ� 7FL �.*���;�f6��5�4�I
�#_�S
<��c���K���1�Tg�	i�tR����p�칤��`3�����ɯ_K����3�=�w'��R�Fk�O.���Л�e}� J�/z۰i��crX�=����F`M��1��5W�
������91�x����b1�&��nK�3�eR4
��ӳ�q��p�����Z�Z�lg��&L��F��l�Ǆ�z��5����MZ�$��u`�G�Ev�-��+1��s�޷�=o�/S?����p���OW���(ibYf��n���xv"
^�~�6x�,V�=:;ǻx�87�=��n��V���dne��ɠ%����(]꧐���G}|x�v]�܊[�@t�� �E��G�l�Cm�6l�\�ӌ
㯝��߲b��
�$���Q�����r�z..ˍ3�R����H�ZL$;�rs���WDQ���j<��Qα{��vD���f䮩��$�.�D����\gK���ǣ^;�׼�a?���:��ed���*�%�������(&Rt�+������z���O�yx�\t��S[�GS�����#w���F�O}��݊�J7�%����X{�3ǒ�a���<�cS���3?�GO��y&��	�
�z�v.V��a�z$4j����$�	V����Q��Z���\quFG�٢��w�]L�D� �����y��e3�lv�# @ƧY9��2��2i��z�ğ��Vn��+	c3"NO�5G�w]�V��E(k�m�r��P�O��A@Г��!�,�Ϗ�S�b�=P���(d��f|c�K|��t�^.kވ]��cK[���1��ݽx'�.+�a-������$e�fxӿ�����B]�T��b�u�-���y�Y���3/6�86�?���?Q�FY���3�M��N���<d����п�T�����Oܝ)Ȧ�%�{v�l>����q�$����\���(\�Ys8V��� �D��Lr�M�Ȼ�:ϭ��z4����qh�دy��~-QT%:z�-�MZ�@-������,�*7��nzЈIarR8���K�2,++!:�܀�CeE+�?کI,ns����\F��Py�o�۵@X_����%p�(�p��N��qb�Z^m|��Ϩ�B��J��'p�P�ɪ묥���ׂ2TnH��u��t4Km͌��R�+p�����Կ?��7_Uݓ��	{�J�&m�W��K�{�c�$�
`H_d*��0�s�x�%#`GeMp���b�ʅ������+3�|�\�O��"�r�%#�����bx6�"d��p
�ar�[������==O�>���Y��1@W�O�ԛ�&�K�|����Բ�>v��	���������ݨ�פr�ܙή������ǋ�]��	q/�_��Ɏ���7,��!������z9؅L��'��;0��ZĹ�-T sw�]�}=���b��{�k�é�xm�v3ͭ7Q|��,���^�_�{/�=:|��� j'���*��=W��d�꽥+�+%^
>�͔��a�b����}�ۡ�ҵ����"&�������Ŏj��0�ˍ��J^r�O�;�pE� ���Տ�N�w���U�S�gp�)��ϐ.���4d��Q����s��]CÅ=�O>kF>������ڨ�'O���3�bN�ѵ �v¥�~�j�����(���ӫWߎ%ޚ���8�9qlz�!4�3��y�ɉ�Am�K�ԛ�}�\t�\e��Y^u��#����O�!y��/}���Fʬo6�����h#�M���;�\R9,�����E�����;fM!�u���o���J<�]����1Q+)�x��AB��?^�����!DF�Q���s)j����o#agZ⡙��*L�8C��a�H�3,�@o��~O@t~@u�jW���U�����-�����	T�7#}]�EY�h��;Q�.-�~�h�۸���/!����SPK�̨����F��u^�҅&U����r��Hr(ܕ����f�`�s�@7���3|�t�����
���/��\�do���ٕ��1��.,�1��7�������Q �egU�P��ʒ��Q�S�L_�<����M�%�F���%z�q���9����o͸�؇�h�uy��
9�>,��Hw,��S��8�δ~x�����Z��'R�1�Y���c���l�S��C�i�C|K��p!�t#�ߒ�2�U���/�4���ߗ�ie�1�����:��S�.�^�or��EW-��~�sM3���:��t����v�G#��74/��jݙ5�ҕ���C���"#���|[��Rv�M������Lu �f&�
	�d���g�eR��t�An�b���un���Jz����&����=���t�tYy���sB��Z�II�\",�����c.���&չT2
�y�OO�Nm��aBX��q_�<��G�yx��
:�Ȟ7�J�ܸl������&Mɍ�C��|�XNx��#r�+=�&�9�����RS(_�.]u�D��N��4�"����#ل�:��΁��kt��V
9I��P��n+��7Cr{r���o_��{k�M��w_�@K3z��;܉�J1�o�p��{���(+v���_~n)�h����$��p�Wc>�}�d�oN�%�]������4���S>0�H�D�-�jל�[�x��"�CaN	�q����'��9g����<�֖���p�P��ZAQ���U�i���9���XE��J�+��&z�H�E�����w� V�+T��dϖ����Nl������&n���_��W�A�	�?!5"�г�`L�)>�y5|5��g��-@����kj.���V��0���� (��\���5��7��w9��n'�,���0ڧ���(B_ �|����I��۱��s��w���)>B�}�ZtK�`�_��ʬ��6����2����2�J.,?6?/#�؞��>��ݚ�\5 md-��ߢč* �@�M�.r�C����`���XY�(����s��-�9}����=�A[��6��0����QL�3��b�o�3�(��_��"�:dJ٨��n^�$�?��!cPW����D-=���,�q8��VN�	�/Gľ,��\c4��������N��uN��m�؈��d�dn���M,���b�m8�w.��Kg�1�Ƿ�������;�{���b���_�������L�R?Ңv�C&�I?yK�9�T��|/'}ǽw��ߐ��13��u7�>u�d�Q�=��7M��h��-����jߎISk�I
6l�Z�����Aᄾ7Ws�!�뒎�p͸��$��\޾`��>��_n��>eU���	,�ѨTB(��J�9�v�L]���0�r4׳Ԅ�S�WiE2ڼg�#�w��PY�K��l���gZ�=-M���3��E�7��c����n�)
��IʵJ�7�Q]{p*ft�삧�'��$& ��R����q��Pm��Dʛ�>�/@���&@�,Y��J�,�V�~����R��,YH=]O���R�bҌ|9�['�lߎ��z+^����zq<%��Z*���zO`�mߗ�6��G;�l�-�ƿoO\��Ν���~�@�o�J4�h��	��*	_��7{�ydvᙉ(�H�f8��zz�,�����)�h+*����D(�}|�O= ���_�xԉK��^�m��oz���f �Z\i{�M\��x�
�"���$� ~�m$�ǟ�=R�������֦�����N�����˜�Ǫ31I���3����k�W �>a�(�ܯ��4���no�|���� ��A����J���@����8�窿��T��*5�0�k�5�닓��^?�+s�1�%Tjazn�`:�C�Kf�O9z�I��*�?�R����?W�+.]�ˍ���D��w���P�'kL��w�2����]Ւ��%��R}���.o����}0|��*'�P��*�0�y��g��WY'��9)?.�����5�'y�יm܏KG�t��vyy9�mV����&�[o�0@�r|ޏ��^��V�E_����'zBW�]Gt_�w��Hްi<%s�S���6S̹�8�3��l�����;o�B}�7���l˵��{�M�gXZ,����{H�[�)�[V���@�cip�9���7����1�[�)�����h�{s�kK]eO���˽��^�t��Rz���\�A�E�nQ%������ɣ��$|��QS�_�r���r����:�ݭ�Cȫ�7�������g�P���
��rZ�33�bxT���iӶ�����
QW���;$�������q���DI�&8�o�n鉡F�ς�j1-���Z� ��7ţ�:9I�JL\���q�*x��-Q5�H ����{�ܘ��%b��_���DJ�SO]�jd�5���0DKw8��Y�e�!��fиDD�r�,�Da���Fԅ�/����Zr����z�.���]_��I��o�xS����¼2�F,�~9i���b�4E���V�gv�X�a�I�אJ�C��wi�m[��vJؼ��	��x,Ǥ�^��A�/�6)�^�u:�ű|AB����n���iӠ1�Xa�k����a��.�fNqF�o��^��?Sn���
��\n�%�܈C�@�fp8�� �V�8���m�l�� _(HH�H��R�Ҥ�WJgmm-�2`�����>jz��v��o:���_��k�~ʺw훽��gH���|�.����AR}fX�,�,�7PS|�p�@�Y�x��}��ē] �\�V]/!��xD�˒&���@�8	Ԁ��_sݳ�cv��f3S���[;�$�����^!�h���4\�78�����\0π�XO�����i����KR����8��脗̰�È#��<=٧����N7�̾^ ���Dp� ��p�b��� �^���V�������j�v������o��ԙR��J'��{>3���suU�tM#5�I�̹ܿ�o#6��f���f�[Z[g�+�� ���H�9���z��.A[>r?������v�Tb)a�K��:�`"j���I=��"&^�Q=�y�V��++'�t<��+��u�)�\X�qf��Es:�Y�q�{b��L4�n���F�'�h�� �$)�|�i˙�3����$�*8��/	�m��������Z���ɇ?��c��q�\�����;�S�G�C���5T�u��`b�i���h�m���5�peŝ=���[������Y/QDho������fg�Ż�j���	ِzj�N� �~�]�j-�`V��$���
�پU�o(�꟨��V�2����cjm�{���D���;E$�(��˰_�#<�%%���@�`0eeev�b��	�
>oQB���Q(4��A�(-�u�� ��H�����uuu7��	�9��IRsuuQ�J�7;=���k�����vƑ
�s�kc��v��F�d�(�3@ټ�_��0O݃*��=.��cg-NA��G��,M�n?[>�XNH��et�drF�Q���ٸ)��M*��D���6�㰬��� ��W��VOR���~I;V��r���,�8� �'�ڰ���~�Y��ol��Lg����q�
;FA�ON	8^��*�C��~�#�镍>����ůu5�\{d�-��s���p�tG�Z$�1���3�{�Ω?7�u����f�E�;+�|��9o��_��KikS5m�a�
&�Ծ�Ӱ�u���#��5e���D6i�V)Q��K������z]ԇy�@K_���O}�:A�pz�
[����~v�Ѽ�����$'K�kF��4Ң�%�S��8�h�$靯�dq�xC�7 ��o��8�т�Ƭ"��n�D�93 �u(�t���d��ʓ�T�n�{�o�震ө�������I��Jt���8�6��|@O�q�q���
����/A}����а�cN��{�m���C@qH+�h5���U�Ͻ�mQ��ge��P�햣�a�ޙO�i���:�[�S�����=F� խʔ���~9��+�}����i�6�q=�:C���-�NϬ̤�H�Kz~�AZI��s�tҳ�X`,�p���u�l���u��:�J.w�k�{?� Yz* $���"U��?�H�l+tȼ�{I/^�H�.���|�=bT��ՄrtC#åay�������n*J������1x	CzL�c���)����~: ��CK~1��fxb- Z�P6[�VPO/1!a"V���2��&5	�[���ttQ�(����ʏ�"���[չ�<ak��)'�/7#��:/*�ՋO�;�J��{k,%���_��;��&���C�7:w:,ײ��,y]tz���;.䳸��w���}���-�!�͞�Ul^?O��C]ɽٵ� 䱄n��D9���)Ig�SĜ�ڦQ�ib�K���o4�d���j:���>����C��`���Sϓ[ZZ�T�x�@���'V�����J(�I�k���)Q�S"�����p��ɒW��b��������)p.,!���u5q���W[lǤ�Z�ѕ7�*��T��J���ͭ����!��ŉ�y���|����*��,�]�y��UR���� N��i��z��r�	��d�k)�l�v�	�RYr<)����#7�����>�Bc|�V�B(<0�M�����5���~G�d�@�%�h�6	Z4��p=��M��ߣX���9i"K�%�ENm���eH�O����I�n�zí�Ǐ$�]�����J�e����_��,���94�H~��.B���k�[�D2-ׄ��8 �j!�o���$0t������~�[S,D����m�zo%)ʚ����ܝ�}��[3��n��骷ز���@#i�Yt��E7�+���~\\<��u~�f<{]����Qp~���V��zw���P�+P�\��(//?�����d)����-�, ����,��\]��c�1uBg��}SO�'�����hF��P<˛!��3�S�Ų�O��qBt�O�*}����̜&�$Q�&�Ukx��j�ʹ/7��';���w�Eꊥ � ���L��0[(4a��/���Dmꔋ�>��_OZ�)�$P��ꤔ��0�¿Y�8�d���������Z�o,_	W�U����M�y 	�FH@p�$Xw�m5׿4
��Y�YKK	sZ��5B+���&Jm��q� ����J5�C���2^ũs�?��.�Z�.������YU*���9^��
>�8b�:[v�x,�\a�|�1��p�������w�x	�_���=a���2x�m/ϓ���І�N����{�:�z~�B�7��ݑ���?%�À+�[��L��ܻw��֐�<�����r��W_���+��G;*�R�`.�9�mN�w��vأN0��/d���i8 ��H)շ��6�/����j?�*s�����)�?�o��!�b���a�ˤ�.��bM��m5�������%���s�p����T�r`�i|�3�l�}���u����S��W+-3�=��tN<<��������Ԕ���Y8��A�Kg�(8�v`��X��87s=ͷ���TJ��,p�t!�ك_��F��������ҭ����ߟ�����U�g��7{*��|���=��d�R��hH[��������?#䓓|�sx����f7����Pi $��or̿~C��F���v4�F��chƄ��HK2��viS<���y��g)$�f��7CqU����\2Ђ�ŰN�k�`��\I<��%E����v9��G�ׯJ��|�ه^y.��d���n�$ ��ں~kI���R|��G�x�����
x01�F�b؟�%��?;����?WW�S
ǘ
��?U+��3�������	���/(E�ė��~�:����S�j�P8tB��VKT��`u�k����R	�%��a���� 礊�N{�	�Z1��ᖑ(j�o8�OvV�+��P����U���Dg-^�����ƺ�uW5D� ��O�kmXv=����ǚ��-m�ʪX��f7=S�jz��L�K�dy�����B���U�mArS �YY@����Llm+�GX������s��^V�؋�>&R�5ꏥ�h����� z{�PU�q�a刽�C���;������߹5��_�U6��c�Hh鉡0�Y�8��N��6Ѡk�.d�/M����R��J�B�q�׶�������&��($|�g����y`_5+N�ț�s�2����2�e�=t=z^4O����bB��lwtuu�;��~�`~_�S|Ҟ0�*�a$�gi���鸤t�U�q��.S�9Z�{6�,�������'�?���9��%B��q}\r��ddO�V#�E��� J��A������{� ��p�铄 �9�k^g�LD�����jGzI��^���ʀ&6�[�����=~�ީ�
��W�W��SB��g�e�qfR��G��Ȟ����YՇ���UAqG�	q����T*i�<:x��r�0�@`�Ra�Kg�_NV��)\��j�����<]m�y�:�N��S�M�|�A����ĭ,��t2L;%�p�q�=��``
�xJ�9䜒̅ݙFҍ��W�t�z=�|tA���|�K����Il�'Lm�)���ϸ�F�0�|�.�{*�_D��b�t,���Q��c�B��_r4p:|;	F�$�ܬ��I����M�az���Us= ��"I�ܺ����K�����.�.�Θ����(�F5�����F|�_XE�!���� Bj��Й@AdS֐MЇ�(k�Q@��D���S�߷����%�ˁ6+Hg\��q�g�9S\�s`	��<^�")"XE�^,Y�<�q�Z��.p�=�ř�fg-m�$x`�٩�~�( ���љ���L�5M^���49��yP�=U��Ȃ�{���>�'�F�9�L�r{��P9�i�v��S��\��[��i�R�/�Z+�xGP��[�K��,j`��������ݚ�Z�V�Or�K5�}���]�*��<�O`F��f&��`���M_[d�C	~���J�/�H޾~�^=c�#�-�ܶ��Ҽ��,��9O����<F]���2)�4�J��֜"����ӵ=��-ǲ�]%Is�����H�ӎ�;Ȱ
'3�+N뗨iiQ鴾������q�X��A�YY�LMO�l6����ZCHo­���(A��w�,������F�c�>���y���e�5v���ֽ�^�����
�g0��{�`v�#D䏏�\k�^Z���v{��Aԗ���x&w��|�_�\�;��f��.�k������/�4h�3�^F(�$��3�FA���!��f�$�O}�/�Zd�b%�0n��M������p�ں:E.m)�z����30@y�P�)�RN���2����Vx�_��أ����SNQ��7���q�.�����=�Y�ev�\�oTR1�'��F}��Bd�7	��xĻ�*׼	�{��=Nv����z���k�������e����5��(�;u����K�(B�
%2�,Ƨ�i���'��	k��<AFH�Zwc���'/X�i��@$kh�������~xI���2��%���'��/j(>��)�.+/
h��2�Ww�0L`�d��K�W���Kg7K�kF���O��q<Q�*�w�6)D�k����Eo{��A��u\�>~���%|M6�@�"��R��[gVsk���T�����ܲuq$\~t@�
e|�3�m�6e$���WO�&��Oᣅ�kr���u{$G�p�����۴1��14"�4�K︌kt�VWl/��R���L�F_aǜ4�Uq%�U�����kC�����+�>F�~v��镉S'QWD$�9_f�Q����t��_B_��5�s��� ��q7S���hW���^��hdn0{g�.���Q1t���hIq�� ��	
)��l�H���������y�{��N�T}y<����R���d)KHc	�X�o2v��:3��,�Ȗ%R(��ml�m4�"�5�$R��;���|��_x�<�r�gι���uݏ&V�!9�l�/P�j�(�@ ,��-���?��:'��ߢ�7���:({�e'����k���۳1u�͙҂�R�^+J6{� ��V����s�k�1\z��=~�A������c7�����E<�$��Ũ%grr]��!����lҁ_t�D����2Tm�� Ut�^�4�X����ݘǤ�]B=���~�jk��`��Q��dx�F �: $�yf���Z��n�45)���W��>4�#�XSyMY��O��+K�A<�{�zdm&�����e@� y����0�ˮ�=pAO�nQRb��!�}����D��Ȭ|��n��,�X�n����U-U�FZ\�%6vvy��r����¥�c>5��>^��!���3�@���������v��X����V�3d7�H���2C������G�9��UK튤���x?g�}|�1hz+o����(s����L?������2щ
ꙥ��>8Xݒ���U����}q������z��0�_���l�>ܚr.���X��=���JɅ$���;�!�I'dW�ѱn�M߭��{�W���Vp}�cNѹ�2l}�N�΃���͜Q�^�	�=�{��r�g�z�k�����j���Iw��	�N�������:Yw2@�^�M!�=�l��`�t����)�����b�ș����)��caU����l* �{t�~��I賕Ҙ1o1�/&"�UUG��tu�ė�����'r���8=�~ ��|d�~wW^&K��Y�D�]�1Q��1E�*�)�� �Ѽ���V�?Ӡ�W{nk�ȗ�&=�K#2��j���]���|)�,U�C�r����!9���0�y��r�]��$�(^c�Y`�0��7��-3o�K��bn���o���7�o1�4o�Ɯ�L����l��zyl��������W\x7B�d˟�:n!�e���@;�0�و�T)��zh�ё�헣7eVRЬ�b���W�����ͪ��ȏ��J�����Sp���4��ND���cz��y���� JĢ�SW +Ұ"�VD����>�"��T�y֪��g���J8c�`f��B�ףt����KB�Y�)z}-T�M�6���_�����%��>��(뛇3���ʛ����P�SoSP�<������R,-EzG#�ݻ��1��[��1e
��	��Rf ������K� ��n2%��@Uh�m�_ �-�؀�K]���Q{���xz�xL�г�� �Y���.~C��i��؄�6�O'��5鿛^�,�Mg�{[u�����Ϙ�1o����ܯt����a�f,����1�t�3�8	m�P����.��|
��#
�go�����+$���5׃g3'��g~G|߱��c�%�"����j��ʀ��S�L����L���A��"�����ࣣ�3.���{��=���%�	
��9$��Y�^�}�+=,���ڍV�?w�]�h�s,�%� ^=:��!���+Wk�4|��Y P��<���"m��Of`��>��ϭ��F�#�����#)�z�usr�HfT<�F�R��W<�1��뚬l:��T���x�怗�J���S�W�}��"9U�o�?�f6^��0��!RG�G���$Q;R��}�r�<��|�Q5r�]Pe#DH�G9{�O�)4��,���s���A	�u��D�O1R	���O"O�X�J�T���d���w
��0g�7���n����ӺX��g�w����|�A�`�t�ܪ���od����6�������.���g'	*H�/a������UL�ߝ4SH��kҠ&�
�$���^��v�Ì��e��ǖ��_�#5�ݙ5��_��.��`����θ{W ���4�(٧�L��ViE�th�����_���� }'��S��wS��9a���������������cY̿��I�2��El~ܩ��g:�"ى*1�\t�:zT��K�ɠ�����ހ���6����9��;�d���e/��5݀�rj�eu!w@:\9���tњ������շs�_Y����24;�����6z�Q�k���>68h�Ȼ��ƨ-,�#~D�{���ϺP����)0��N	7���Lqe���+jrr�:!|g�|��;#��j/Z�$zI�u���Sd�Gd\�an�&�/
�m�|�`Q<x��瘸M�ٝ 3m���lNFV1�N��n��R�S��Ɛ>_0C� *�NQ��J.�H��J-n)��x�B7]�4���[�O�t���#Bs tOɁD���xIS��&vO���;V��-ώqE��YL}�
�U����(:�<;��O%wa���G�	�lAU���x�ɳ��U,�C��d���i����%�5qQ��>H&ѣ��0H�W�����::H�⩆���pGK\�
^���G-g|.���5�]�`��lUK�p޿ױ�m��p�U�_޿�mow+�ͬ��3C���������T�+���b�c�(<��sC�}<���CQx��އ�c�1?�d�(!�nR.���Ŧ�\���&��i��&M�\����,ӎ��M�2+�T�����}��n`��ؒ~��*����
���c*�#)�չ2�1)�$z�����p:��3F)8�Q >]��2�皛���@�A�9�A���Ìd׈B�>c�c~Ӭ�ev�������ֻ������iт���Rl�;.]�Sz@5�s>�h��A��C���O\8�])Ma�"�	Ji�ů_��uB�LMNF�`z��i�M�����`���v��Yw����h�σ�̰R:�-	��z��\�2_-0��W 5L%/JsG��AQT#��>��Ǽ��)?r3�9�䝐����z���?e���h�/ d�wJ1b)�׏��҄���5=A&rrB&F��;y�U�c��\<�>���WO���-~ԙ�y��v �o�V�� �ŝ�4��>:��D�/8׏0��T�(�<�D	��V��B.���sun��8b>������E'�����E&}�>%�6ؕd� ��\^�Ǯj=5O�����=A��&�P�D{�;����I���)�Wv��� E��sݾ�L2��]s���T��#QA�w@����~Ij...��ښj�?~�<���'T��K��/������ c������x|�7������^^��rqV=�>�f�v��-�s�yJ��ߖa_�(/�4�����ky����]x�����K��W� ���?AX�vab���ˋ�j�LZ�6���"�וkL4�=D$H���+��ͱKxN��	�|d��(�p墻�o�)�vY��ZyC�_�N�<41_;�?Rx?��8�Ae���O�K���i�w���:��P�$c����5́��4[O�3�^�v�¨-FT���:�/�|��-]�q*�n@���?�S��7� ���xYm��!��9�W��m��&�w�x�ѝ��)}0"8y%k�����9��#x�<Kcqj]��Uu��۱�ýi�m�d�Ӟ?��l)�����	�&j�RN*%vܵu�~e�ߢx�=��=0��ۅ"mY	���7�]x��>$�0���^(}u�Fz��E�F��G_��b�<�%]�EF��|W�v�#0H�d�ŜhL���s�m
�ԓ4����H������@���pj��3�q��he}�,O��P[¹3�J�Ji-���B��[��6:sҏiWv9T���e�H����)�����hr��w%S0�a�퐿��䴪�y�d�p8�IxIb���J��f�92�ܠ^d���~$:�O5�itQ�i��~.?8�a$�V�9 U+x,}Iͭ�̆���<�f�>*�V�1���.�m��y<�f��K�����M�^m���'ʗ��e.Wu���[��\�ߕ��S��XK]h^���<F�Ң�^J�/i`�Օ�J9kACTT��2���R��|	L��M��idDO��H��VCcl���)dX�I6|:`�Y��x����x��Lcpu�MےL�at����gMVm���R�ג��u�F0�k�j׸��>��} � �@f�&2V�a���E��GD���8�T����`�Z�}��'9��� ���U�)ck@�s�:��͇{����ȅ�ia��@� ���-��(4	����q�����2��V��W�{�����b���{BAJR�I��#�=,w���s�[��2������E��z�6}��$یd�=��a��V�k=������~vm�_�>	6�țp�tx��=�Q��؛qg�I�]@bջ�������n���փ�(�E^͕�������LV�|,M)�4���r�92�C�!������"mCG��Y�[�){�)�.�2����b9��!����� ��t۰�j Q-��޾;���{+���M"������P놛,��jp�\�����/���N|.i�fȅ���O1��O����t��bo��p@�USW��3|�;'Uģ�����PΩd��cg����L�d�woa�u��$�'��k�b�
��;
G3 IU�W	9�m*Pm��YJ��Q�XH	5����\f�������A���"R�j�#������o��-�#k�EԌ-iK�߄����ܮU�t���},N'�ٳ��܂��B�@c�j�S$��٥���[c��@��1\"Y֭^|;�r�C2�9�3o%r:�q�C��Gq�/�JܞWIU�� l�S�]�yv�o�#E��"&]�?㷁	qY?�q�Q4W�J�qŷ�x��Z7?�x�'[�	�%�c����tF��R��N�����f>�N+�M��N;�;5�n' ��r��7/���EJĝ/]�߲Cpl���|T���:���^��(0�"�2��C[;�t�^���\���yn�,�󗘝Ǘ]>C�pz/��tr���	T'�������b�T!�\L�yzI}	�9~��c=<��k���5v��JF�9(����+>7���Mk壣���q��O
�H��FGES	aÜ���e���&kI&�"@�= �X�"e�)3���򗹅?��D� 0�?D��:���ʨ�J��H�t�������tb
1�1�bk����<���&�L>�v��=�@1����X�I�Ն�_��۝獫�E#8&˗T�{'��A��?{m�{�k�l��5M����;K��sh�U��9<C7Y�iz�����䭭�����{��pD��������M�<˔���W�3QY�T�1WI�y���r]8�'�0���).�B��SM�%�JY�E��?'������-��>�y�K����R���!V=��a1�C���)�[dhp5I��k�z�PcC����k�:�/��y�2'�T��Y�O��9��ԺY[�N�����"�j=�|@�	�V�g~�E��5�O��^��Z��Yt��)L���Hȴ����$����x����]��\T�Ǝ-ѧ��%]�2���,_ꘚʹ���s��Z�Ai��nX�t�~?,�������=${��^���L&3x���0N��	����:n1�<�����~	"�N�6�
�n���V��2�4Zԃ��m��`��R=�r���X�%�_p�y�&�
��"b�}���'� ��Sb��@'p�!��̲#���4������w����s�~\�?���(�������u��;zu�ꛊc���<*Ty���)R0	%��â�w���s@��t�� �V�A��t	F�/��ۂw<��F�m7����E3��ջ��^��� �^�h��ꃚ�M+����=��şt�JA)���G��`��J�v��Y�Bz�Y���"��|j��'�A\Wڻ���Y�%l�C���տ%���i�R�T�?��JB=��Gq� ��� 6&xEN�c4���m��������ѤT����#�>�����=w��]'W���JL|1�1���@>�^=����Q9������`�X�Q:7�9�D�c0��xg�Ջ���"�y��k���7��!?�Ћ��X⳸w*�8#*Xz� �b���t�/1GD\؇s�q3Dn}n8NG~z+=L�;��_!���������D	''!�*�{��[Y�[�j������l�L0�~{��;���YQ��Nz����9��n:��/0�*
%}x�>������`sWܞ����({>`�)h啰���"+G�O8dę�X����|�^D���y>�iɏ�r��S���P~J� ��(���Xw�h�������M���I�;6'���O��]���P���Z<�Jm�:�,�y��t��alb��9�rD����=d�-c(� ��2��3�H��
 M��ySJ�b�;".a��P�ቀ������قq��z�-�E�I�r�A�I�^H}f����f^�&j��~K�u��R��|6���sُ
�4�����2�?G ��ypaY�r����}}����h�s�?5b ��?��M�ܭ"�(�t1�[^����/9�o	b�\�'�,���Tc&˃Ԧ�}s���!A{K�7l}'���0��TV�z�Pq�"%\��َ���~ђ:�%
(��g�*��㦽7�5�Ɇ!������Z��Ů��[��Gd����<��ԯ,�9U�⬁�ֹ��wݐ�k�?��?���0�p�ZnM���=�w��9� � `ޥ����ru<_�ŉ>b��}#��s'>X��PT�_����]�V=��76�>��H��tr���<���}��Rl{�8t���P/��!���/_p���j���ܲe㑫O�L&w��d�~0�o�$#�YA���{mӹ��|�6��~ޫU��!��)�����ME���Y&�
'h{�m:��T�����4-��?���Ǻ7f��	��UF���^�\7n��g�6�ȯ����"!?�	Kټ���v����--e�Լm9��W��Aj�&����Cj���Q~�._��3�S2.F���B�A��@Y�WWWuO��p��U��\����'�r����q[��u�\�y��D�}�wGpNo�2��viga[���c޳��]sW�<���#|a��ˮI��a���C�����)n�]�K�yk"�td�].�myֿ��w�!b�0#P����ׯ��^�x����mM���-y��T�_�ۺA�I�;�q<L4����[�E����#ù5�@𩐽�hf7^�������^?�LRg��yyjy��� I�{*C���^��_�?ǡK�6~����<^�+� �����-��Q���>Ai󬻻{���?�^p�>?A�a%�� �����qҰ�f��H0�EH��-I��G��Ə&�n�]p�6�B���ݒ����'P��Hq���-������ܞ���o��M�����a�7�wG�ߥ^���4ܸ[T�7�E�e:��)
�n���	�B�"K� \��ZZV�~��g� i
`;��C޺k�OvRh���-��ɬ�9��A�C_��E��������U�-��j�;�J����	޹�T��� �1��?C��ِZǰ/�
�S��r��Ĩ��fؕ�A�y��B衭���iҼ	.4
խ�sZ����uJ�M�$���M�C��mk#�����z���8-K�c�(�_.0j���$@�k!�S�i!�ID�C�TQz����-}���AD��뜀�	u�/�ݛ!?>]�������� ���1�?�7�3�NÛF�X ��3�\߭�騞����g\ذ=��M��෉d���@����O�p�S�_c*�D ���k�J%����Fa5-*���	�2���y�/��<���]���`����w�N8o+״?j�U0���c�J����0�{c�L�[״���~!�M�X�s���������P�ftil��w��3���v�����%� "7�HBiM$�#��U�Y�̥�SPr�1��OR�?m��蹡��2s���(.ew�m�珀�g��:�I�"�����K�>ӿY��~혓��96���+�����w5]>ɧ�
l,Ӯ� @���p`6�����e��y�-�"��Õ�S�)�U3�It1d:Ư�)Q5OҺ2�c͏d�� ?άh�� �?K:�{�GD��~\�����<X���4�W�V���mzr,٠�x��9s��po��x,����Y�(��ۭ,\\\_����(�S,��W��TzuF�J5^�:���R�q�B���lZ��5���-٫QP�Q%�V����\Z�-�/�x�?$��Ĉ�1M�y}c{.A�ņ%����VY\��Sr%�5��ap�/�����Q������7�J��}�A�B�%����f\$��2є;�X���1?פg9wfO�2�~y����J��u$$���D�qѱ23]����iI�TH����WGXN�����ٳ�8�J��3o?M�_~��Re~�����_�8/0P'\���NOZi�����~���ÚCӞ�9���̕K�w��n~M��Ir��ks�J����vD��DU?�PJ�}��rr��oC?n���d{��\WWWG��˨�/����L{��?�5j�t,�I6��t�M�G�u��c�� a�qb�^"���Z瀏VU��O��7�u�}z�9Ϋ���ڲ���5�2�USݸNRVZ��ę�)v�}���-��\V��~�1�@��J�����m+MC z~}w(�!�z�A�dΎcAi���4�3��/跾6"s�֘&�"[6��ͷ$0�#A~zt}k#�����,��
,���FQ�o,�|��~�=��E �(HS�O�;xQ�;&� H��Rf����n$69�S�W�����,5�xA�}(�3�J���i��Y{���������@��TnIѣ�M߻������%�L��U��Cn�r�щلS#2 ��K�t?t��xb��Z�zn��*:�ߋj���%5��O�zv�?�L"D��s�1v�Br��|�V���<�[W;�$��fh6b�t
� ��n)ބ7���^^�SQ�$0�Ѥ�Xfc|IV�6�w�ךX�Sc|���-7��FQ�����$�?�OS8P������:�qސVчsr��יc�$��n�۟�x�����h�$p���%�Sm`�����p\�I�{��X��-K֐F>���L~�v��F:P�H��'�KG���S���j�|Cr��^��!<6ᖥ)�*��(�8b�2�K�˩﯇�l�W����Y�û��џ��r� �~4�HkpŏEql=�U!#_�t��DY "}O��G�QW�P׾�/��_d\$��n=b�������·�z��2�6xLv�q��c'�p��}h� �URW	� �L�g�}�r���h��k���i@�2��`�}���4߾!Cr�1�l^��&J�7��znz%-	�D.��|�P�@�������t�P�dv�����oV�GƱ�٨�|u"�n�j}b�Bu�}~#p�K��jm���ϣp�v��8��H-H���!OS�Wx�u��\s)���\� ���|	 o����	�^k��KF�@���6q�D-�$��eZ'P���ӽ�oN���wl�y�cTi!:=�̻����'�)T?�S��UZ���_=�i@m����C1�Ā[�o��j��zB87�y� o���8@� �N��f��/:��� p-#���ԕ�A=&r ���^��a�h��ى��>}\6`Ջ�3��T�ѧ#o���Lb��t�m��s��a��>��!"�����푂j��!$��8b���R4Go���Xd���>ˑlMȾH%y^-������PB��]�4�v�M>]�r;�[N��
��D
�_�/����8V�GIdR�_�����_i��z1�����Sj�)�d9m��g�uK	@����i����O԰8���/m��}pAfN]�D2���`�<3��0s�'����D�W�]O��=愯��P�y��B���=���9�
J��8'���_?\�d�lD�n�>�s�6X��V�(:~/йa��Fz<��E!gD�-l4"��K�^<"&��a6�Ń+֜�yC1`o�>�X�A��eR��� �����X.�DQ�'/�\!ї�lT�Ձ�t�����2�����3��,�!��n�7������z9�ІR.#2��M������T_�O������/T�>zҾ�ԛ��O1K鉳�/�K�:���epJ���}fQ�}r:����'��C��]S$�b�L�k�v	H310����x�j�k0�������Ŝ:�j� u�!��8g^��I���޸�#���=�L����]J���>ռ��A�}��'Y�x�}����2�j��vLV�f�>r�Y;�@	X��v�����*�;�7��pQ���8x����A����@�����z�m58�b�(&���/���#���)��R�bN��W���GΙLh�!�Y�dG����J>��Y�>(��Q`�lB7�o�@(�c�I2]E�����i���Ѫ��� y�j��ެokY���� #��g*�I�w���!����c��G���̏�;4o�U������ߖ7�%T��$2�)s.��iV �2�	�U�X�ڽ�s&%�ycw��
�٦�����)N����",`���Y� ���Ç0��O���`BbziX' �O-���s�r�z@^��I(�}�b�Y�{������Z��n;������������Q�@��u�jލ��S3��k$�|f7��O�N�ԬA6E**�@�L��y��[����H���r��v;�%44�u�����*J�9Ar�k��� 1��50��4D��:�5EC9�? yVd�������󰼏�攂����Y���q#?��t�yTzX��}��Q ���w��5(�(��פq1�>0�Cz�A�@m*z-�4Y���M۾�;!;Ae��w���+�a~
T�\�>}Pt�/g��m���xlE�õ'z}�/�������/辧���~�m��?WWW�ތ�m�w_SS�Z}
�� ��,�!e�h	[Y[[���q�'�NGӿ��+� ykop����K'�-��/B�g��Gį��?�4���[|g�K6Hk��+��R�vw/��IU��T��󪯍��7�,�?8h5��x~@X%;���:���E��f���E�ˁ��g�i�A.�������;6�m^�3��j!�պ�;0M��h��<�Ա$���|>������Z��am�y�i�:���<�m'���g�P�D���� Ô���olj�A0�H����)��q�c����Q\O�T��y��"�-�q�ыb�e�!�����+.��Mp�q�~Ȱq�D���� Iz.lؑ��u��O7����?��"!~�i�d|���PD��+7�=�C?ޛVN�2�y��sڋ5��:{�s\?�v���hF�?��ņ�� {�o�#;�RDy<�T[~^"�'���D�����m�'�d�_�0�-w,�_�
��t͡Ob���ԇ��%��mT�y'�T�vBxr9��o��x1�rD$���Q�|�^r������YxX5/q��L�mw��gd��{�[�)+���:�K����m�� �{g-h���#�jt��&y�G#�Fr8z�OH]��%���&��{&/��5"y�n!zU�
�4������l�e���kt�F�a(����^��]���X'�F�"������zg��ϑ���¶� ;0�i ���l��7������B�ut�xj��|��Z�ri~�Tw�q�ȴl�?����B����ﳱG:�<u�KWr��w6��L�eu�4� ��Ų����F^���-+01�J���
��%�o���(N��7M��U�&�v�D��˷�J!z2Y�d^L���O��5�ہII�!m
9���_,��&S�J9,�R����U��<��`���gb���D���r)�_[S����t��)�\��N�i�to�>�\	��+���@���L�uJ�r=C��2%�M���GB�}Z����ON	+E8���5^���|����N�*ec�ôLW<���xu?����s\����_B[t���K'{2���-N]�opSc�&Q�whk����bg>��O��V�o�.�K5��ߘo��Gq�$�Z�g;_T�@�;:^'�'��.O�B[�
Lr�pЅ7,W�f�K��w�.N�!!!���y|�i�:��0~��x�4'E�-��=�]�j���c�����?��,��%B=����#��&�7H��D�,��S|�Esu��<����]i:���#L�n�Â�c����֛�Ė�P���ٮ���L�>
L�M�ypAb�\�zO�����_��y���o�E�趎�`�R����;�M+�c����e`8�k�C�Y^���bb����fy_��Euê�f˭�fD�ڵ�`NN8-���̱^G6M���RH���<<�&�ߺ�9R+�p���x���r~RRRR+@�=o{��{��&#Q
|#�p�������A'��2�T�����L���"�dN/�>�Mk�-�K"��F�9��>}m*YjC��y�ɱ�)G���%V��ǚo|��Q��M�4���3��q�_��9+)��$7��QRJ������}�I����JGTX _^PJ������#k�Xy&�BJm�x��LJ�	m��,t�Ud��,�����ʘ�-$ե��ñp���g'/�:sh_���Dr��T��3�"._�HF]��y�.�����r~S)F����2dv�E��jǫ��xyӒ��R+3�h�:���B��Uz3�,����MŘ��ϓ�-��������%�����8B�h�e�G�(��GFFJZ���
�U��e�g��L��x���y��Gޑ�AW�˷K>��kQ���FN6�ˆ橉	��Poy�b��e�=�rg�*Js���J�6��U�7���ie8$29?lM��ȧ~�T����3�
Wn�%Rs���l�WbҔ��f��?ۓ�p?����5tJ�����et]��k�R��b�?�b0Sm `�K�n���������f]%��ײVb���� ���Ã~�8Jq��<R��ݤ��Dy���@ҕt�~���GQ�h���u��@}���k���::Tg -�'�RA�-�$���s��f�|I~�K�k�*�iz�S�{�j�������݃��BN�ܫ�AEh�?�z|��un��� ݣ�l�V��ǈ�I&9�<�և'1�gKn�.a_�����P�f8���;!�V�bűtBBB/hB��O�r;���%k٘������#Jma�� �e������B˜��&Lb�?o!��9��"_�3���a4Ddr�K��I���~�V�㮿_�i2��d��D�j��`�QD"����WUj-�a,��<��r��o�Q�k[�e�ӗHN"�Q4?ɸ�썃��Y�i�톈�F���������k��_�~w߭2ǭ�J\���V�'�7����3yj�I����0�*�ɬ������BA��,Qo�01cCfm]���4g'P{�a�+Lj�Ru&���.U�mԢM�:T��^�[`���?�;ȴ��:��A�b.�}�*=pn潜����>Y %J�Vy��/jr\�?i?C���:��20Ni���$-�Ǚ@T%�AEU��i����{�Q*���{4:%ؒ.����l��T���J�����)|��(������O2�y?0/�آ���n8o��*Af�	?R�h1>�K]��9�zE��A`�_���==I����
��F�h\s��F�Z�h᥆[,ʐ�����2d�8���1����M���@���I�"~oO^q<�P�x>���&���^�]U?R)x�Ƶ,l�Cj��� ��k�N3D_El��"j~�+Hq���1�mh��}@����V6�M*c�Uy�u����R��nȵ������{~]�+���5ȏէ���K�z0HT��$��Gq��.VV�Q���}<? �|�_C�/����@��^���I����v�X�<���UsL\.d�{��kC�l*���q,�+�rsM��Y�?�,)��V��iщ#i�Z�m:c�c�V����7��,�7�v��Y�)�3D۹��i}����	����H��Hk�9�}i�q��[}�ij��p6�"����m,�~��E�2t���Mq �8��<�'#�Q%�0:x=�����V�Q)6�I�u�g�l#r?|�`�g=�:uAS'w_��vH�KRp"�p�˰���=JxD`;`rɆ6|�%|,��fd�[�:�0mHDrE�v#��$Ve�l0������ڇ���r��pR:�I��1�2�Gb�7���uaaB+�Y�L�o\����91a5�{�%w�ӛ�鄙���ܠz�4'�;H�̑�T�	��\X�I�e)��8���2�w�,/��tk��A�<�B#�\�q����5�T�`�@w1��2�qJ�����`q�_[G�O~V�$0V�w�/Ps�h���[C��v�X�o(�Mj�HP�
��]ё�G�o\_�R1���i��0��Q�	���%��kf��9L\\5���a��K�e�!� ���m��s�ꛁ�'�Q��q1D��9,���F�{kz��
�>�2��F��a�
���%��009�� !�j��ݱ�a���q�\
�Qy+1=��2V����:�X���ku�-�hizf�n�m�#~� ����YEf���&^���
�J�˪����/9SD�M�'��������᜘�_g���J����j�ۇ����_Ә���N�\�K2قT�iE$M�����-���g5^�F}CՏ=�'ċ�A��ƨkW[�4[��HF-���B�|R1l��\�e�p��>���v���gY�iD���4qfRU�LP��}A���l�A}�`�����c����UL�NCZ��aKs̕0�s%�.�2�`0�[,����&��>��\Ú�M#_�m�Q=K�9]zrUY�����T��(�CX�=ڃ ���d�W�	�(##��p��z�I��N��:=�1��h �(E$����ɩ�V�O?��&f�U��"++R�`�jȯ⊂e���V�� �t�AL3�F6ra��0��"��ԧ��-~(>����99IY�z�
V/|��J�k̈́:��S���ܧ[����5��~͌=/�aPf�P�M�Mb--e��B�ߊ��5P�r]��e����N�l�hW��,�7�8$��r+���𦢸�������D�01\2戮4�)�|&�r_à+$�2v�E�_�#f.�x�F�E��o��P����^�1�d`���DGv�]ܽT�
�Ó	���ބ�1���@R6�j��^~}��CPP��m|E��$�֥Qe�:�)1����g�A�2	˾τ��E 7<��{~�K�W�-ş=���4�[�RPZ����1%�"RuFx>�$t����ۂ�aX,��?> �**�"��^��Ҡ�=��5�k�?�2���^jm9gT��[�ك�,\��e���ќ6�C�L���NH�g�;�G����A����|H
�6��_�2���1Bh���0�WXu�?�t��2��Qf/\�n�%�� U��Q�BJ��`Fm*� ˿���bP��w��S�Yݛ`&����Fu;��sjD�X����z\�:vu��|N0�1mucj��C�q�����u,�m	ም�^~v]޽sl�>�v�/���y�=J0�q+E�s�(�}w5�;��=�c�G����������(-ً�
�;mV���
��.�٩Gk� ����@I_��<�i�4	��uT���"�E�p�0��}R� ��u?�L.�|�L���n��J�%�yD��	g�����W���%�m)��$M�ʓ�n;��?ئ)q�5��+���P�Y�kb���J�,���׼�&�{�m����;~cKnx�J~��-�*���#��\��>�:�f0M֫Y(Y�;ϲ9����d����#lu��kO�+��r~i�^��0� Q�V2y��4ۓ��ia����T��yok}ߦ%l����"�n�g��n��k:~�dQ6�u�Ifa�3��)9�! �l��Ԋw��f%����cэ�pgp���}����֊i���iCkRb�@�uN�w�"J�-���hi�����z�+�֢�5\v��IE�ņO9[�\��g��Ζq����r!����$ɠ�|��';��������������B��K�܊�6!�Җ�IJ�/W4'/��� '2Q�\e�ַNN�!������U�'����i�Qͻz�Ŧ������v����4\�a]��ק̘^aN�Ou�����ڨ=ja�?��}�������+N7/����XD[4$Ǫ�}�c�Ȋt>�1�o̖L�g�m���Ee��I��Di/�`�jx�S��4�B7b?�C���h$�E��6� ��N��@�-:�ӀH1��:���f
�7+j��Q�h�Y��TwR��5��L��99�����?i �&)/��arE�נ�X�ts�4H�a�U�&b�N�~�5O�`5�\��(�_&׬\,נ\���� d�Y���Q�����9�O�H����_�z6����o�ˤG��9:C[�'W��dV#=��ӯ�D ���.���(~% �ly��]/I-�z�K�����$��rs�i5Zȅ
>�._�N�<��驕��sz#Q`�eť�[;x0;k?�XU6�F�X4��=�\��X��To��.F��뱊�:�a���s��$T���3
��ZG�2`�sXW33�bf�5E"�Rk�?�˕;C�^2�j*��{g�����\��rr>$x��� ���8J5:�/����17�gW1@���5�Cz]��x�y�l_��ޅ��e�hw�?��bA�7�{�,�
 i:[B��x+������@��>��xl�N��;k�d���]i���,<����3��������Oެ�;��x�T�F���)���x	N[�eQ�{�w������Hr��\|�Ԛɿ��1j��F���f��k��[.'ʽ��1;PP�nRj	&}��S	I�!�cIk����t�+;*P�`,�}=��(�u��A�Nz�촫ꋮ���c�'d�NrW�\w�{;��U9v\�+�$6	�N���Ym���	�B<7�(�}�aj#2�2��4���e5C�\����"������)ݚF� C��~i"z)��q��]�����F3�t�� �SV g!,t����Z�[�Aտ�ӽ�����c?@Z,�I�����,�B��Y��,o�'"�u�l��;��n�?č�ٜ������'NH�X�eՙ�׼L;�e��v4j����1
.�AޗbB8�3�||���C<gA9U���;��2ۭ�'����y��N�=�p�Ev��os9�{U�8��m��	��Gz��=z��^��1I�!�ar渚�.�߂bI�9ڋ;!6�*k���Bu6���n�`�M�$#�i5v���}a���������:%��e��?ܭ">h�!����S��H0�#-��LL	��h�������l�}���5��ef�vC�0Et7�C}|��{� Λ��J���4��[�@�y�ˠ���"��#���TT���r��=�������x(��Mʞ�H!�0!$c��lI��d��c�����al��oٷ�uEBCv�dK����}����'3c<����9�u�u�	�4�z�#K�V;�Ahեn�t��w��+Y~~���b��������Snc#�����/B�ܿ;�Gu~�D�PVXtJh�]�Ƙ���v���ތԴ/:&F��$�U���I�ŹEEf$*�Ȉ��b�RE�X�0�7+Ы[��� hݱ�,�'�_h��4�I���tfv�����$;���67ֈe�~nKz\A��m�gq�V����V\���?��)z��g��\-�?f����p�G�_~8u;ф�E#�.
�j5j���{��g��gYߓY��t���5�!��� ��{s����p����$�+F�l�)K�N�̳	,	s�_j��v^���/���� J�Ϫ׺/�U4�"��$t>h(�����.��6j����m��d��� K�� �2��̚��|��I)3e�􅩝��+q�o�|�-d��x3Vh�=voubS�;R$دnOK��2�LQ]S�5A��ϒɯ<�8翙>�(#*�#
���]��k�S��9�BI:�VW_�n�뽠����㴻�TL��t=��.	�'0^ý�ɫ�0��-cǴ��ƭ��=)�x��s٠��h��7B���n>^#�&�n�?U���GI-Tv!  �jJ��wǔ`6A��T�{��k�rq4'�����4�]��[1��{�M�J;�;5������D//Y�"fS<9a��Iܪ�<k�&_���y`�{/$!�=�T<ax�x<�:��v���zW_R��̣m�/ �X����%�'�`��I^�-�G�+.(��v��k�)ذY���ʰa��ǚ�3k*e���J1[4a��BA���l�2���}�g^�x|��k�D��PFd�UhXm���*�dO�ش����7C�"*�	�.GP+����k؏�Rg�y�,j�{�^�����g�P�B�nT�8��kۤNhOQv��ء�@v�N$��=�B�g!`T2�^����9���~ں��I����ډi��F0�̊����=;�S�w�^PB���7�ӯ]G%�&k޾�m��4E��IX�����/.r$�[(�����D5oBp�k�,Cۈ�f7�G�1s�����EɨHA��������!�w�Q���E���0C���jX������	����z<�	g��rA����B1��3,��m7i�`�X����-�̖����O��/{yr�-"3��z2��r~Ө�}3�B擿�>#E����d=����������"Q1���y�|{J*�D���рW�ֺ;.A���hT�nZQ��<깄��� ��K]��mEi��lP�\99��u��`�o�v����Lo��O��Y��K¨� �c*���z���T��:��d�+�e�,�py��h�%�{:���۟���B�3�d��g�����s�vWPm^t�2��n����J������T`�;&|�^��m�^q��f>3aB!���ԛ��-N)6Ƣ

��˔�>��Me%��~>CVè#�Q�̦P����e%��0�<.�jȻ��w=���m�h@ͦ�f%��{^9�IW��;gg��D�t�z%��B���w
w��f�%"�7�Qϋ�r���,������-�^5�_5'%��R��P�'x
�D����/ڠb�֌*�y����[[�w_�%�{��9�
&'�r�i'ѱ'�i����]{��%���(���;˨�L'��˦5Ų�I�q�6m�I�ѹ�����>=~��5Vs����oA�M�P>A�(���|��3k���1�WJt�Ӆ���l��jtP|���ZTt'Ug�`�8-K:f᾽=�%�;�z��f��N����W⋢�������t�V���W���G5�ʼ�O��5�H��rTZ�=���AU����s�x�l����$�80P��Ԟ�)EM]y�eqC�nunQ
J��ys�J0��y��x`���e8�~9���Q����hxLuRE�%�]��+�������X�,��E������fz⸝R[�e`����|�'?&�ӳ��6���,>���
/<�p�A������K��ʏ��D�$F�������������yէ�`��mO��g�d��os-5� N��4���/+����"�6<��fk�Ʋ��Ǽh���e^�8�y�i`{�RO�����hP�{��U��Vv�:nA����<�B��^(+x��Lг��!�G���W�.ېs���7�բo>~�8�������O�BP��0��;�
4eOVᄷ�j�-��p�Ohɤ���/M
Ui��ŒݓS<2����{�mg��T�-m?Æ��UC��8kl@��7V0���v7�k���ג����Zs�8��Zw�&7Mf��57|��LY�k��捤��=A��1���L�:!I�󨉂��5�JMgkgGv�2l�a/���[��~w�0f���W�` jq�5b���A��\�&�)vy���f�([z#����)S��lV	T��sMƯ�NY���k/ �ah�n.n����}�	%pV��h��&N�]���+4�l�Ɇ`�y	��Z�&��)�O'#�������	�V�y����+��t���3&�����v���p�������>Ē.ߛ~�Y,a��?�ĒU۹2aߎ��蕛�&(X�Z�L��IU��>�/�e���H��e`Zz��\_Y��	 �;�(���@u�ߧ_����k[3v)�ZW�_e�!��鸍|8=����S�Ƈ��2C�V�>h!��S��u�����ü{=8��Q+գ�/�}�PA>�ꣵEV�Z������%#�IG�=u�������dU�'��d��;�7� o�P7��65�љN^�:)�w�B�ŋr
��**\Eї���K����yH�4z07ː��=�{��2S{��<O֠�����W��rq☩��IsR��U����p (�=$lﰽ���$K�;��ו6˧j��T�UX
^sz@�I���b�q��#�S�=�^���mgk�����\�!/��ۿC8R����	��/1B�ZYY��7`��\��S5IXDboh�� {��鶞r��[K�տ�`W��k�Q�<��4{Gڎg�:[�����]}jFZ��e��W}��A]�J��PM�9���${���`��	��hWl�Y��u�w��e�b��'5+싡'kߛ����[V�?ι�z�
��s}D��Ӧx�h�,Nj=]��VI�bb<9C��m������!�n�/n�R�;T�^yj�>#
���z�#^��Y���D��F�H?�j���9���1%
͆`�#:�:$]\��Z�d��;�1tJ o+f�ٸ�a���P��|G��r��c� ��������g�3��酔{��K`a/0�f�N�Fff�0�[_*�Θ�eD���\T[��I�Z�����nX7G�*8��Yb`���Ғ�2L���a�8 ������Ҥ�r"؃C�hKY�K�D0l�]����3��*L.��7Y�9|����~D_���7�]�g�%�$δ7��62�Cr��Z[��M{5�Om�4��Kǯ��eM�2�%�Zp�^��� ��Ï�<��[�4ɱ���-���i�	O �|���i��6�ɫ�Ey��Ѣ�����VN`*�+��5����5^e�u�Ǥ����R�Kw��?�)Ľ�g�|�4��f�\9:�\q��NI�z��	*J�3~kGP8�,��V�8J^C{�G8TE^K�B����z������m��He���I}�{x��P�a�JQ�n�D���ԑ7�h�%��d�8�t?���z�S��[�mo�����9��{x�BXy�2�z6���*
�JHHxԂ7ZW��d `�c��:�W��g�>��i��C��	�<��Y�$��)�8�b	��Pa�MD��-+y.����i$�JL��#���4mBeMC�H��'5��G�$����Ɯ��?S�������[cJ2ȈP%N��x��Hׇ�8�a	CR|�%l�:�:r����]ra���FaW���^{��@�:�%��#?������j�s	��,ȞC�s�aF�|$�1���&����_���N��Υ3�mmm�)�_������JTR��=v��LAǔ%��C��ݓ�k+� Q/H�:���G�n��ܕ�N^:�P����ܬp6x<��)��ӧOi�����R���-�H�	�C��I� ��*Q���PF��x��P�,�g>���*�I�n�A�Ւ �~TQ��������˒�Q��W�n�kF���c�\c�y\�^��Y���N���6��g������/�;�$K�A�p��E#�7�x����4��W/i���r�^Fy.n̲9]RU�+�c������S�")I
+�RIDZ�~}oơ��s/�,��V��$��� �-nF<�<7�*�&�/ٍ�}y̯�/6��@�Z#�BU���l�lb`�K�(]���E+_����w^��lL/�����g�5�����
�.O�MS�y��]�Z��ͯ5\�����!��b\e.u�#ЎpWXC��@��J��i�� ��?�5�01-��K=\A{1ܰuo$3D��?p��=Fw�؈%�E���s_&Դ�k��k9x�%��(�x�[� ؐ��Z�5/,bu�Ă�x��M�Њ5���O���Tg������}~����@�=���Wj$+�m���ޢ?9���)�4�%�*kX���{H����'s�Q����v�E867���<}ݟ!�ۋ��қ�'d��GJJM,5�GV���BSt���;gOD�&!�y��R�0"��P�1���i�n�*,��;��/�c~B��L�N���{�%	��Wt�A�e�i�ԑ��ډ��i�����̿�\�u�'?���C�$�tqFZ<�vXt����s�p]��8����B�ߊ�]�������`@CM0IWp�Ǹ���G��=3
�E��'6��l��.i��탗�l AO�s�1��X&^qHN�w�;rsKJ&&�o-�����#D��߿ed�[W*t`:�v?L&�5�/�٧��:��7��l����,D����U�%"��V�/c�SSS��F�[���N�5��W}`�~�2Gi�c��p���LA�,��<�3^�<ۇCů��aS�sS��K\-䅡����9/:�s�b�EC�|40�||�Zj��]a��]|��{�P���x���s_u�Ƈ���(F���/��+Ӆ�x��4w����E�����S���+���
�Jj��!��:�[���?�}��ՏŶw�� ��M\uѝFqIX��̠8B$���-��ƍ-=H�$�+��O.�N�`fCeT��`�x�ƶ�ԯ�P��J��1�'؀�J�I�g�"L,���99�9�n�4�ح����!���Z=�d1���;����$�7���U�)�|.N�.]���O��u�me�m�88�W9����c�U�x>m'ժgO����O~6�a�%��p����ӪJ���<�#$�ϥ$�����&=���w�=͍LLd�m�q���G����N�zE�}��J�f�h�
'�[����&%�N�vo�Duީ�����o�ߨq59f��� �'����H��<�gS��*���#^�ߛ|�Y�="��J��CJ*��r����N���,{TghKG��C$�`g��c�1����Pe�{������������r��D � _{<��*Y��7��Xy���M���-�SaJ�`�pC'3~��
`Wϋ�-1MF�;2	&�c�Q�,q���q� 0���HWַ�oV~X�/4^X��~��. �[�J��̈́oH�o�@����,p�d~�6�xw,�#������P�!����>c1�_�"G<���~��ob���HC ��wk�\L6wk���JJ,{������(�W}��~XGxĜ�,�<ʌok�D�q�#�u=k�Jo�#le(LV���F~m��N;We���R,�bµ-&���>�X�I�W��b���>�;�H�t�Uћ/օ��P�8� �m��&�m�����\qA�z�]F�{n4h ��O�Ozjbз�Q� �Z��y�Փ��"'��و�j��Ӵ� ��r�e�7��&b �p�t�+���i�����M���:E����s)��ΥWQ�N�������˞����
̙<�沺��`�a�]���:.�XD��vǢ���Ew���{��l�p���d?�{�K;���=́!g�T�M�/�/��{d�+Gg
�hyX}�<���;���<��~~M|�E#�H�xX	'��������6��Z�s/��JCW����BFx�v�ăl��Ċ�>�����#߯*��A�H���Y;���s����݃h}5�VT�A�K�p�ܦ�w�a����&�����h���鍁�ӻ��2��G�UP"�6���٭�q�s>�bh4\9��v�J9Ӧ��_ˑѰ����G>�*���.dz#�zn5@�J2aLkm�0[p���5��[S�@�����z-�8�2��.���]5����7Oqw�懓$3z���z�3Ur���Z ͦ�����;D��t��ܾ};*[��xXF�Y՗�����a2��>�5��"{�4�gʲ*+�H��;���_k��?\�-~y�A6-q���|���y���.8k%w��'B�#�2S�`�j���ŭ�hT=�7Q�7������eUOX�6��7�~\k�_�N�4�N���XS�^��l�����s�� �Cv�(�4��K�]VB��a�?��ʟ��<}���p���l��i�뛋��
�]bK�3�Wc�>|�:t��\^~������m�p�v���4�R���}^�)��)5:Le���,Q�J�3��=�f�� ��0���p׃�,�վ���nS�MU������&��TN��0i�嶂��m���ֈ�-���/�b��qOn`�N$���>���w����޼�$��]cϯ_��
������ju���3�bb��O_딶���bT~I 	�=#��|U�]V����g�|4K����ܺ�R����Ur5�*���ܜV�eAS�
��5&&�}l���Ob�4D�>$��偡�c��N @������<��V��z����];O����'}!GgV�fͣ4�%A;�%aAK�d���ᗽ֡E�s߅�"��&gB�NZջ�NtB/5--����3��(�Y���Ͻx�N�q���&|ML�ě7o��mvL
�[kN):E��0��>*qZs�W;�����dm�̈7�r9�����Sm/Pn/$�ٓwW~�9��u�����(��v��-$�?0i�l���䯉����owz��
�PR��_���'n�i�jr�rZn�&X�	 �L���PਐoBOe�m�����>���j���^��Jf,	ra!�݂3Df�N+}5�~_#����X�������}h՛7e�� \,1�m�i��	��8mr���<E�����ݾ21�l/����������Q�9��k]�'xG�����J�Qϙ/w�*�������B$���i��.��H�w\��H'U��u ȫ��y��_0��Gk�%�@5��̛���B�ɽ+���<Lտ����w*X��&���ϗ~M62ǰ"����ѡ
��o�1�p�;�v<�Zq�AƐ��5�ܷ���7�N�d>�$����%��&M֩�j�|����Sm�9���jlEg�h N*�u!����xdAҺ�)�4JCC�F��kg٪MN;T��/0i�{��+-_�d�.@�/��s)׬��?�ֱ�!����&��W�1sA6�A'�26���u�c�����%�G:b�to��Z�R(a-�Y��-��	(�`�
yKK��������ۍ�"�����J�&g�^�x���;D9�1��q�7�UY��'G%����G��J�e>�)�8zC������f�Piʰ�ZZ%��ԑ��&��[J�՜n(��K���8��b�Hy�1��<�5!"X�c�P*�rX#A�v�Uf&i����[߭�E�ߍ8<"�q8�G~x��'_+�����:��Q���9�ɲ#�t6pm%$�0�e#��@,K�G��Go*�(�h"�r��t�Q%�2���z]&ɼ��8�Ckwg>�,�X=�m��;G��S��¯���g}cՔ�S@C+�0�i a�;�"�}���5�(�էh��Ѝ7)�t�������``f�3s������ޫSO��S��1b��X��n�պ\�l��9������L.�!�)��-�a8��6ZP����N��i"n�x��e�?�7��rI����H���h�zމ�W~����ow ��1�b|vr3�%�^���+k��W+���&5���]�������Kx#w`Lzu̴UV%�7)�C�/�-��e���Q���lwJ5���߿�I��a����C9�^��f��t��M��K��.���K��ƿ�������gatU+�Z�k�)�K�L3��Q�J#�\�C��@a}�)����V�ky.����m�����V̄k������A�����黺�L�:T��.�� ���օ�|�Y^���Ц��Id<��祜O&�0e.D-h�yV��La1�#��qj	]1�y*fԕ3�0^�[N�f�N��w��<e��V�yۻϗe�ֽ������ ���˰	�ē��/������z��� ў/Ǘ����m����L�
R@U�T����D"���h���)7D��ᩫT����r��q�΄5��́����
�_��MUR��z�f�{�?C`���Ps�������}�}C:�*�QU�w��w��#6��*�9��g�-8%�2P�8���LS���D���p[ܥ��	7�����14� <P�/�)������i�t0�4!�}��*YLµ���!)�nR��vŜY94Z�P����>�7�?9�	�S�C�jF]��4:���bGU��?��3�s'n���^�vT��h���8EM��%}�M1�� ���V�V!kV��o�py5%���Ѽ��jy���"B'�	'z�ʌo��V�`���PBv�gi�W�E��.�u,}���M��ʇi_�~hikSj]R}��J�[��*lJ��\Mq�#ߒ���I����
�yV���'�g�P��%�����*1�WQ�bHG��?��eb�O��(~q�/,.��k����%l��Ύ��M�}�z��#:����͡&��˭��Dtdz�eX1611���~[���������T�ݷ��x&:����Ϯ6)�#������M���-C��qg���Z
AV�!���+���i0���F�s��}UC���
I�R'�g*�j�:M�w�k��������Q���,����6e��먹w[[Y}m���dzXgg�����k:'��r�������ẗ́�'+e>�^k1T����A}+�O��0*�E&����ܻkT�l�v|F%�|�������H��UX��&��i�@��jO���X��E��LήC��8̣��8��ז�*����i	cj��Ԩ�|��7��cZW��Q�|'�e��������cQ7��T=����p9�������Y�+JR�pUT�m�[�ɷ�±����(l����;���yE���G�a�g�W	��(�J
*���6��7v��R�Z�Ǩ{"�� �j�67�c�:����żS��#���}���9�!*]��/w��:��:C\��"�ޤ�T���3=�}�4����ѯ���5$DP'�{�N�T�u�8Ai�TL�b= ����
sR4�����M��ϡ'?���|��?j>�k�0����nNpS�����DH�bٞ@����Űɘ�'����2�x���k�\���o|���V�x���H��F�>>>~��mx�TTT�Q�lFUE�a��� ����p�Qr�Wk&L�Se��#���&��k�Ȓ��`p���
��|�wc��G���T��p�>�O��,�a�P����;��\BB!�$�"N7���5�z%���b�gP��=�n�Ĳ#2"�Q�0�3����o���˛�6`����c��}Ht�Ć<X`�E���0$v���Gd�sIK6�����j����!<�������Ω���JD��F��^X9�E}��x̉$w�7�������w�Ps�FP��x�-G2����3pQ�^t?S32���ʱ�R=�Y�ׅ�����Q��"��S茐�)$[r%��談�ڧe�����{�Gzp���i�IO�ҏ�\r�����8�_z�Y����3�× ��3@�-�R. h����)#"hhj��pcg�zR olV�1��-r�Ӱu�q���B�1�v��[#D;���כ9tE�r���l,ʌjf~�V3+���A�=��yT4��ѡ���~�gΎ6뉪�G
2��4�[���_���Y�G��b`z��l�i(�=\��?��j���s���u���h\�UB��8�Q5��
�>�}��Q 
�g���1UaE�=�W�hN!&�$���T�<oG���Q��iu���I�2�>4��,Zt�'镳P?�X�h�h���Ee�hr"�_Ư�����]�閙�Ow�5��q0���b��K�z��x]��2��H�-n��#@uK�]d��b5 �6X��Xtkdv���N��� ��k���L��E��¢��Ƶ�t�ij���v�%����h�ԗö́�j·��������䁢�7����� oW ^��w�@����2]���%"#�;x$G��9ұ���J���,�@����:�ô�����U���|�Zd��c2L%bQ��E���h�:�Yꙉ��E�>�3f�+S���e�z3�a���#^���2=�-e���%dz~����Ml��sl1S\�x�x*΍��G9�Z�0{��t
�\�tp�_������������ ��هN�{�4l,Ȉ�a�E��������X`��[�nܸ�A��S$���z|&�i��8K��"�T�$�)��0O��	����Jsވ���(����:ޙ[OY��o����J���;�����b�|���'�,z.�񜩚�==jÒ��bɆؑ2�O,,!<]��3r��eM3I�N8�7���&V]k��r�%��Pp8�&����p��g�&f�g5X[*�Q�%��*�ee ����M��)ӣ~f�k��J\q�&��J9DvX�0{�09ejf��8?��x4�f���Oț�r���/8"��)��=�_M�$�;�F��f�o�R�G�Llן���D����±���Աܨ4##�N��}<6C+���L	il��='*)�7�z2@DO��n�%8�[�+��BO�H%k������ Q�g��2,�<�$i7,!`G�[������V줪��eL_O#F������5����:/��}��oy���3I�� ����ݛ�`��n��+ԧO��\�a�T��}�^���3���󸚰��۶Ww���'=Ha�73��j����%NOe�`ܯ�z�caٰ\&e4U�|�	�h
�����\t��`�;u��n��|9`+���gT�.m��&!q���[(a��v�|��%xMZ����3J9t�\q�$tߪ߼LZ��ÜlX�͍u�%��dl�\C��ݙRV����b�-����#_1�����b.���,�YU�i���7�o�����>�o_z���H�А�V���_z�����#%��=⃲[{��@�	�'/���j_���If{kpJ�|���X����!�4���f؟��u�������t�a���/���n���;����9��H��T�6�6I�:D?xN^%�<��CO��5�>ZW��,x�j�@OPG0��T�Qq����l�$�a�t6"�./�N�uT�d��F��=80 h)�v8�ȏ�,E�5�j۰��0>�"�+�!�;2(��:��6^Ev��z��H<�hf�e ���>I)_w�Z������V厧n����U�k�X��b�\W�.��I��z�_N*����A�yAD���I�h�AQ	��4!�w�4yZ~ۅ����22�:"h��쌙�;� �d�ib#J����bȻ��A*��޽���c�.��	K~� ?v	y�iM��
!a8H���H�bB�C���;���}pd'�u錿��vQ�He.xh1ɗ�#m:��1+k~4*��v|�b�����B���]�A������ݻw�ZkMk��d�o?�b�:����g�������g��N��l�9Y�ѣ�X��b���5��Y4\�J~lFJ��
G!�Q�+� �!�m�����dQ4B��Z�¹
�,oE�+V�o�>Pea�"*//��,���s�|�ġ��X� �<�P���t8'e�~u�0#�R�&q�Ԩg^n��q��W�����O����10 t���9wdVb���smJo�g1c}=<�/���{�#�`�z�@`��7���E��Έ��ݺ�u�'��5�}[;;ã��]�x���yPl ���A7Y0G�$�2Ip���}���x�_��~}5G���}����-�Ͼ�"���íQT�a��c��ֽ�w9r��.]����I��;�RM������p���pb�O,������IR��].����7f@�<��ې�VE&�(!������E,�DG�i� ������/���S�Jw����H6�����x� >L(�n�]�8~N�XZ�/�^eG��7�iB�c��¬� ����|{3o?V�j�z�@b"�Iae5y����5GY��hFE��ϔ��n����-o�'�w�;e��˼ɠ�9�]��.i����zw�����<F��N�/��@4�@+[�v�/�]�@�"�:VL�)Ho�d��y	m��:��ѥ��O��)�`�,ƈ�/������]y���T��6T�vL��-p��:Y��=�d���l�]��d(��_!>�k��^�E�;3p}�/����G�,�GHCSަL�#�WZ���L��������b-�����00]��7�i^��''�a}(�n��˦�Q��xmBD�K�!��+��XMj�K�Y��A;d\,���Mq$�,��v��V����պ�~9�X�rẻ�g6�/�Y�:�r��t�W�Oj�#��)���|�ɵ����a�3���y�1��hbd�Z@�u^��k�O�,p��g��b� Ogo�X��~�%l3�Z"�DR����Ԥdq|j�f%��S'�n��{1����t,s�ö�<&�kx9�ݢk�+.�8A,쇓��y�0���ς�c��<X��g\1���ɩ�xa�V�_�����e������?�V��;[e�O4맃���*
D��`S��(��kUa4�*��k?2 ���~���4�5��=>M��m܀�vX��0��{��XB둠D߂�0EL�j���	w�����'�~�V�1�����p��Ta��A;ט���M1�9��T�T�]�����K����|1x��z(mv(r~��+@��ƪ�y�ECr����[4Ԝ��M�x�|պ݅���mpPe;�9:A��,�x�8r����/q��~n�-'���ٯ�Py�d�ng8�Ql��r��c�_�� �*�Z��ޏX�;C�tN*�J��)ꎇ~T���-���ۧ� �u-I�,|�������z�¼Uܰ%�9'�NOP]�
j^=O��ѥR�qM]�a}-m�/�b�&�d�<X�[L�IZU���ݯ�)s�[�W��.n�(y�jXv{o'y��>A��g"~�ڗ�fq���Ȣk�)fѲ���W���˴���U��?]i�	k=NȠ��}ڠ?���vS��c5��Q��Q�'4�wr}|p��&Źs/`�h��Ѝ>T���CQ9�f��z���ɝ<'�{�u�~G��e��$)�CA�����~�>'���I���BT��8���u��O$y�:`3&��ն�*�R5������m_8�
Nƴ|�0�ϼ]���<Zʭ�~Ik�#Nm��-tge��7�#��t���Ѓ#���ԭO2]�s��S<r5���}���j�Ϩ�B��i*�.�3-�dmڟ��07s�x�^=�H�qf����Vѽ�3�#��o��+��x���gRҾ�^.B�T�@��"����5U�/�4qSL�]�����qZ`��� �ܓ�-&WW��Z�vv��RE��4�+.�l��t@��o�O����ũ��"��2�������S�׳�*������_��>�'ܣ�����Dh�����I$b��x�ҭ�t)4�E�t�$\�7@]�%F �3�q�|�d�ݨ�s��8I��ε��lNhE�m��KnW�8(�;kh6#P�vo��},YnP"����T|����<LI����3}�R��r�A�V��۽�O���x�}��	U:��t�^O���]i8��!��O0,��W�����5����T�}K�ƺ:��ׁ�O1baa],�N�f�y�4��!���VG�W���0��ى�
�%������F�s��w̫��/�`�쳘�� �I#\��d''����f�!]�S
'd��V�m�z��fU�|�qS4pC(i6<h�ﾙ	�I��x2l�	]z��WQ,����V:�҃O�Ǘ#4Ի�X�`
e�~Ex���!T*�Lf/��������˱H]���c�;�+%ړ�� ��/?�MvZԼ�����SH��.�����l�m7��ց%7�ᒚ�XUU���������D�v7�>��В�h�-&xe��A~L�!]	"�9F��ͼ�V���g�#���f*�b� �o���%`3}�����
d����~8��`A�XOlT�M���j/���G;��Q/�I�.[�q�=�0=6z���y��A?�e|~O�����~ܸ�sn|�H��u,_�Y��������F׋�_��O���}O-��hqI�|�B�T�'ۼ��Z�R[��ݳj�7���*GEE����f.sr�ۓ��cb���#������uy���%��YZ�c=�`9��N)(:k�"�
F����E��\vg���+@[�\΢
�؎_Q��kԆ�����y�&��=oa8,�3��'�6��ɏ�h��NuX�gՔ��~��15L�Y@a5WB��4�����c'\�{}�{U�����R���z���T"��f�3G~��JM}
x%�p󟡫JzC����UPw��=�� AiUb�?��Zfh�0uA�oQ��5~�I��D�BK��5����I2$~f���e7��'p6�Ha�2�ߛXf8�7�H�#&���č�b�����E���'��(�g���G
J4�>K��+x-���w���`�!���	�Չ�f�<ݧв\5��]\2�A]���e��s��HkG_��6�Z+���!�����j�2b�0mu��+V�W��"ɨ;���]�?��H���z��L�z<Vs�_#٬��<8�z3��e�Z3�BT��#ܓ�����i8y%H��#����b�~�w����N�����?h�)������r�|�CLi=�e��y�g>�9cغw(ϣ�������WjF�	bɆ�2�"q������=d	�+U���j?�{�5�2�*dj2�ս��5i�o����7�m�i�&iF��mB/�>������
�������^@�M�#
�/)��� OH��-��W�x�F���-�/'VN �eO�eRBZ���y�|M�c݂3��
Oa��Ҳ�֗��N�5�-��Oq��J�~5��pk�F��G�������3Iq��h��su"0��+���z��Td�:����%��t.��q��r��w�џW�*��om��T �M/�\po�&��߫�»JQZ� ��T��6wsgw0������v��ݫ�4�ǣW�����^{�_]�	�������z�*�����.��W��]�<L7��i��Y�?T`����4bl�Ou`HJ�Ĩ���M+N.!��T�-���+w���ј��(�����|�U1B�کa	N�(�z3�����[J$)�1H�×�T����c(F=s̄C��2k��ǔ��{�4�Ov��
�e��3Lchpآ_�8%[t �,m��L���DVU�#m�R�� �{%D�D�fQN8��tD�u�;��BU��uh�N�|�l�Xe3��~I�D9���ȭd{�����<wg�	�TT���xT�/-���WGOA���/;F�U���q�W��gΑ~�ss�>�p����>e���ľ��A`*�������*^�K�\�9��(�B��-�����r�+=ܲ�}�>C,/��]�����?��e?}I���3Ń��.��=���A,�7Y/��>^W��ARvS~
�����i�C~�rsq@����Ħ�ĀɦM0G�w�Q6����=6��̩��+WZ�����t1�M��<�C�ŷo&�g#/=',8@�.;��ۇ*qB�{xxx7�X�Nv��b9�q�5�2�ӡ��+�w0b޷�5j��\�����}���u�eH�TE$�Y&
b�;��8����+3,#<�ݵ��:���{���E�ɀo�E܊�<4��hćc�R���f;�q�ami銬0�Hp>��=��������֤�I�l��Ř4LrNIIɏ���K�u�2����Ca<�Tߴe��j�zύ��d��Y1V�j�z���O��P4�6}	�ܸ�q�����]-=�Z��Jp!ټ��MQ����G�_"��^ Wu/����Ez�V�i��O�Qf������M���C������6����OR�R��+㱦�P\q��&}�-a��*`�6����e�u�[O\����$_����G��F^p�#�:>��#�%f=�x���SdVYII^�1;{���V�a��ǫ�k�2�t��1]��xt�.{�Ut/������A3a�2c0�|�*8���^��I�|��+?���E$Y�^LZ�y`���Zߥؤ6:dF�j����	����7;w�"^�"k]<"���L���z����ej��1)�U�N����4�F$�222~�û�,5%N�Tj�{;�z������R2�4�{-�����kW�&�Wvڙ[D��#'h�}��d�ۃs�V�T��~g�M�y~�Ut|��y1��7��9�C��a�dE�}1jvR&�S�,�ۮk�+��ǰgF__"�"ǭ!4?{lǒǐV��B_R��s��n���z7�M���#�G3.�PKR��ӹ��d���'��G��KG��J�K����t�
=��	��DGq�X)f�k�2�]k�7nX~K�M9�/)q��5}J
�[�)��#zh�^�p�Bp�r~^�1��Z�]k8I��J�m7�
~�o�y�'IU�����=Z�,����̕���]p�p.�������rrr�Ln3aöG��-��z�?�]\�-�hn�1�uw�8� �p\>~��6�p��~�X[|�\�ы�|���
����7w�>%6�z6T�l.U��N��v�24��S-O0���ẅ��6�繥de�fɱ�CZ�N�����'�N<x��t���y�J���^�Ԍ��(/�J��XM,�3p���~m=��/>�F�3�e�I]8<>+�c������ۈ��T:
b;�1����$Z;�Iehk�}��tE˱��u\ؗǲ�����������|R��ڍ6ڀO_6��uΜ���D}�7���q����v<�5�q�����LQE���ж~@��Rގ���s�(�3����g���)�o4�7`,Z[��8�H���o�;�\���h��-K[<^����z]P@T��L�w<���?.�%{����J��SfH�8d�MF��ބ���#;���$�de';|O���w��n�p����u�߯�u]�E�Tm���h�Hz�H��E�6oJAk��T�]}�۷e�d>�2'_�/SE
L��FUWW�����sd�	��b'~eK��N��#�8��% 3y�"��R1�*L�~g����nh��LM����TKPE�cei�r�c�𛼶���B8�L����D\�1���������[�v��q��%C]ݿ��?�i&�TNEA��wޑ{�=e������ ��R�!����0X��wۖp鎝���'�YC���w�l�^P'G���w�L�Ȍ��~��Ҩq?�vv����5�)�K���aY��x����� ��ne��1�5�r�,k$��s2v)V������{�������A�е�f��!}��e��gG�~}X'�b.�0���
�Eg���1ɓ�F<�ž<���	��u��(��?C��N���`��z��r�@�T�-b����~we?��_�Y��=�vB�u�5.I�0��"���UJ�p�zu����B��pW;2vz���	(t���~���=H1������w,,,�qɓ��"�5��Ȉ�1�Y 4����*����:�Y�������z�az�<�g˜$���t���C���P���¸|n�6�q�-5ъ��~��Z��<G/s��6JH�TaVn
�QU�( ���$��X��H�l�w��U���n��2���Q�Utt�4+>��A��Ŧ�s�d��а0A99�����3\�bҗ-�03w��YV�]ݹ¯� T�����7�^�=ުn��z�҈����z�	�.t�-�#��u��'�/��`ӳ%�i���5p���A�p��R\�r�V���}�E�8T�T�MV�!l�w��^�&e��4��߿G&&B�����Z?��	n�i�g�<���x��#�������T��N�j�����K����v��qaʪ_n�^z���Ty��5�S�)z��<$�������'�|!C��P�@3�q羬r@��\�Y�C,�;��ﶈ�̇n��J���G�"��ڏ���M`6X�����3Q��*&"2���ˋr�u���+Z=̦���?�짟���E��"��H*QQѷ�i8�$h�˱Yۻ�:<��g����F�2�����<�bD�=��TT��+�I=�doܜ���֖o��F�FM˷�t�ɱ1��F���݉��*2\�``��q�bn?[��ùPϵ�?�k�e�4�S2�b_�911�0�ӕ�1g�\�'2��Ge3U��B�V{�Z`l]��7b�U�xU�d���1W&�{�:�Jl�Uu2���J�ﳢtx�>PI��Ie�Df�ka�O�㪫��Oֳ1�>c��Q�S���ui)[��:�3�ir��A��7�\��j�H�k���s��RD(�v�7��j	#ht��vWZ,���i�8��C���ى{o�wn�9�՞u�u��s}�0���#~���Y���l��@�9��bf��H,�r���-�B3�r?�7\�����{1�?�M�ߦ9tݢ�����/M��Mjc�@�y�"[`uuuI��Z!w[�A*��)e�x�¢d�`di)ب�^z%XQ7�m֐o�3E�*nF�aBuad�m5�G��VٴD�):.Na\�*�R
^���������s���E��Y��Jq��LT��6��Nf@���vJ�*��b_��������I#����� ��|%hbT��.�����K[LF�矩%�k��eINd?�����k)���>���?\��3��XH���T9���Dr�;;ک7��%�����O�F�M�Aʀd.�ZN���_Z��NF4�`�1X�0��ɲ&!���\�%	ٿV�0C-F�e�ux-l�_��0�ק� �=��8K�T/��kzr��O��)�S��0E�ύ�z�<�ű�LA�P=��|g(����������"��ŷ'Sn�s��Id������=�"�V^��;�̿��\]+.����`�>��9�O�|ja�O0��+Pg�nP�.{:
Y 2�}��`$w�P��h��fW���d�����6Mmtn��?8�ۮ��U��x��(�)���5---.ۖ�8���2f�XJKQ��ϑ��y��G]�������'��,�����)��E:�j=~���Jז��+-m�]��������bA�b>a(F���raw�[E�D�e���߄��9�Q3Pn�o�دk;��Zm ����/���U��G��ueƴ���ܽo�Z�3!�-7��Q�q�ͺ�w��V��吇-[�����á�\�(՝r�Ţ�J0�s��|g!\A�Z1y2�7�Vtx���YMlO�;>��i�95�zQ�ppp8f������%���LL�ם��PB����g|--���i��A����H�U��� 2!�O�h|�5lΉzF���?uS���]N��b2BIP� ��&�L��o`iG���=2;kw|^�p0i�7`z16� cJ'jljZ��?����ۃ�������p�e|3�\9����t��L� ��C8��F���?Ϻ�Q�^�G3N���N�������wt*�Χ�T�zQ/''஋e{E[�R�����(��\MPJ@��Yͣ ?:`����u��iΝ�5��T������[xp�X�M	����vS���<��+�O)p�fx� �ߐ겊������Ҏb	���Õ�|�.=C�Z��7�+���B^�4�djt~��XK���Cώ��4t����\�Y�S�{⌋�\)��TfM�+_eҝ�C��\�v0�u�B(����ZY��F����
�ܗB-:z��B��)scӋ&U�d�ɛ34J��ۈ.�t��uc�W��gfO�mz�	*UO���Ζ���}z�V��w�ϧB�𱧪H�U�i��U�B�78�Ɉ�.;��?uW�}�H�`W�0�߷��q6�.l��Ų)�\���^Z1U�R$��6��USGW,�j�p�j�4����~��������}=u�ޚ���"bb?��?�,�Ժ�6�4#���������Y��ϛ�Ua_G�Г�LC4�n��������Sl�"86[n��ꑤ!�A P3��SEe���ݧEL��bc2�HG^^޵��#�b��l��i�=��5�3_9��/`�5?YNC���Ɇ�P��B�ľ�ee�;R}O-}n��E\D��"�?�w���f%
)��;�@kTU|�a$�@���%چ~�W�Gc���|n�ւQ����]�0��J�8ފ/��Ͱ��w�<��vW�4ͪ�����p����zʨr%YX��p��
�{�N�Yr"��͑����1�B��~F�f϶�?�O���l ���S*��:6���&�禧�a�wQ�)J0�n�m��g�d��<eWV��\:��Cͱ���w�6BxY�F3�a��f�K�(�i��v�ݼ��V[+�Q5��`N�ix��\=��ߠ��m�\����ҧ����=�(�S�(%R��}Դ�繖�t
��8�Q�eL��F��m���L��`�-����и�v�]��b�X*y#�BCCH�x���Y��44�B�|QY���w?����>������� @�F-�3�R����O����R��ZN�9O��Sm�s��Q�`� �	�-��ʽY��C�_ѵ�R������<��2�� �n��7v����ͪN�wxҵ����%��QE��.��	�֋#w�8�"�j*��5�Xf
ٱ|S=���q�����ߔ�~,)����yH�����AN�e���-�P?f�d;��7�����!A�f �B�Bp'85:���M��D�%U��|��N�"����K2^����z����� U!���^�����Ey7x�fW�G[j%�2�Je����$XP�"ԫ�ַ?��0�۲��^�`�j$�Z�9>Ģ��/��v�M�#)����C|�����O�m��»7~���1�ս5$�\y7��խ��YcB�)�e�F}� ��g�[�33s��9>��/�����/(�aggWbL|�D'���
���>˧��7����y�%	�H��*|Z�+���ʊ� s���Xb_UI��6��{��b����`�U=tu�ⷈ��vd���h�=#n�	�q]fE�$�W�ܳ��ބbG�*Yh�_��=|G"��Ǜ�}�>���xU�qX����B���s���v�B�c}�ҲS&6������Ď�Ȱ��@�@X,����*�����͜㻮%�=�JY|�UÓ��B��Xp�͏g<۝_���s��W�9O��yƉ���|iރ�EF���(�I)�� �B��b�(���{-����eW�dh2����"x��<
����dM��Z���>۸Z]ځ��.��e�ۖKY�~\|(K�Y�t"c��E�}8r8D%+�Dn�&zk���ё���/tކ+;;�=�Z�v���æN:`+�1#��� �d�IyS�i|i�����M�r�֝��T��>�T	�K� )k�X����f���u�&�5TQ{t0lCTo�=�A��e(��%����/J�J�\w5Α�t�Fs5����h��֦����"J��<���yVi���]���EHTF/@���ɽ��r�o�&+[�NP��u���/�m�lll`F6�G�/eP��
�J"""is�R�����˜n�\�����+7��!��"��C�qT���mL2Eq�nzK�k1�(մ��Z��0'&&�=;�>���#S�D�x��	*޺�#C�����Qh���Y�듛�{k�<�������Y�T��2�%�q'�+�n�/NTH(I��Cw|��"�
ϑ�sWC(��Yg��>��	��u��N@E���Ի�f��.��>U�(s��*�>C[��mi!�A�,�i�0����6ZP���eb����݋2� Į�Ͻ��w?���d��Gl��
��2(�P�>#�]2Em_~��M[A_�O���G�>Od��mm��X��fN��O� �q�*c۾>�u��]�6f�Y�[j�q�4���1��2��%~���緣��C��<�V�x[����e�.�J�d"޺V�d�j��lzV��E��{�(���%�6�w~�i�0��PZ�z��,��!���c�u���t��&�~6�ٗ|��2T��l�QRn)���\�T��c*%�&�-!�׵Y����I����;��g�sy��Eg���0.Ѽ�v�-?Κ��{��א�[��lCXG�cߥ[��"�2b`�à�J��v�	�u�Jp���
�*����O��^�7��^u�+4=r�����Y[����3�����w[D�N�"��/ɚ<v����(��8������0&o���{�2L�G�Ր�Ϟ�L�ӻ��p��o�.���P�l�隥��^�)�Mo�p�	�j��)��LUy ľ17Ρ�0O�+\� L�gQd�a���}�2��t�yJaX���v7ؿ�3J_����9�]'�>�|w����W��9�,/�F��9"'}۽+Q$� }�:�Rx���5��������c�x�Bw4p9+�/�
n�'�ǐ���𷅫��������``y=���E��r\X �1�Ɩ�3�Z׷�t�\<���y�w��қ���&F��j.���./KM��m��{��h@{����X�:��@���Mt-���z���ݪ�Q����F(A�>@�gZU�_������!��h��E0A�q
�5Jgk�_`�YJ0E��{F�8x$i�ƃ�d��ݨ_��|�]ן`ȗh��B�r�}�<JSn`�5φ8�-�ن�A���}��� ���D�d.FW�M&�_���=%^��0�R�)��44���￱�h���\��CLJz�.fdn�ޛA- �VT����1�Z�漁��� �i�E�4R��o$���E��6�Q=ʂ"eQ���^�P�����ԻJYC�s��)��(�W}!:�O5	�޶��5|�_4�<�<�K���ܩ�;��uus[n���Yw6U��EuYr2�}�L�Z�o+*��N�n5�{" �+�B�G��ۗ�T�c���{���^V�ɕ(���w�LZou���SW��\xJ
���f���>��hhh�{��������a�W�e��0\�M09o�^	FF$IXɠ��fo����� ��[?���t�k!􄲋J�Æ��P3��u�;�}�W=e�%Q���T��G�_�b�	�5��;eD�$r�,V\>n4~r��J�����N���k��ry�3^yU۱��-M������_�"^�'1�}mm‧�j�809~�P������xCq](�y4����p����my>\H�ŧvKݩhv���������.a�闵F����_D�oW%p�&������~�x��g{.'������쟸~&�ny�Ē�5T�֎Rڢ<��gBj�#]5��2�A�BbF�� ��7��G1.2L�Ȃ�%��9��-O�����7e�i��A=j���\��A���Ǜߑ��Ǐ���0�}S�8(/jѦ6�m���P���v�T_m���[��xxŲ\B�[?�V�s�����G����;vr+>� ��,��|p��A��[-Sq��~�e�U��N93�_���uUי�x~~�y��H�n�޲�2˼ʙ�r���8�0'{b����2��<������lH`��ī����=�5��E�5���A���N�^�[eN(�&�t�1�)Wӯb�.1�)Ƃ%$j��k�6��SMc[[���b���������^�`��3Ԑ,N��e.ҟ�y�2�}ޣ���N�l��f��6>�Rpc��4z���Tb6��-��v!�2��f&4�ٓ��U���"@(OrGN7�ܩhږb���lii1�fd`Px��zl�������2�D���	U����@��g_��̟��?��uͧm��E[W�o;=9-Woa�������H� $��,P���0⧣����'���cB8tˬ�p�}�у��^�|9)��2��EP��DĻ֪@uB-FÃ&�<�&�:z�n�z.�ީ.�>�Y�~�ܽZ�
���w(|�#H���'�k������fE�:J����z�CY���uܝ%ᶬ��x9fh���Z�n`E�S&lE;�=����;}u��Rm�����e��*��7qGB�|�(�����}�/�N�~G��V����?�ى{zz����OT5[ES[���s�\R0\a�X"�Ng�ay0Q� ��O�h�Xn�Y�{�e�Xn�48����ZFD�}����]�W�TܔG'�j�k*"���>���bۻ����f����4�깔6��|���L��vN*����M�?�T�J��lZ�fp��ex����O����R��R���d!�_�7ir_
^�}3���t��ฝ�ϐ��8�Eы���W��2�D�b�yy ����4
qV�.-�w��Z�N���U���O�Dޤ�Y�/����3��Ȓ��L\��.�W�xbd4P�� ������s^a�u���G�A�d�0�ŷ�߶ܩ9c4үe�Y oN�Wd�(�]����h� T u �s�s�#�O��_&��u���\ĥ����5�
&	�ϖc����	����#�j/�⌁L��cj�t��܇.٩���P,����Sb�� ��ǐd@�w>]2\c�Q�Pz��Jf&����9B�X�,d���#/}��'�ꍑ���T�2�U�����]"�l���dP�����_�nV�3K���������ϟƻ��!-�F���^��R�J�Gy�uTD�C,@~{�\�~LT3�^P����t���My(t��u�(�M]Q��X���"k�����~�����F֖<j`ڵR�x[���ן��_h�ɲ��)a��[jS�ѿ��Լz�_�����W`![��C�BB	G��=8�����u� ����R\�Պb�U���[\�Aޫ}�`Z�q�6��,�<u�W��q�0 rx��O����T-�e�yN� xT�}}���}���8(})S� Е��e�t�YB��j�U퐎Ŭ\���`0=�d{� ͵5��Z|nVba!���宐��F�k�Xt���{�v��/4�1��?�ܑغ�.�xp˥o��i���s��X;ѣ�'T�5;%�p�@ÜkvГh��ԁ�˺'EMWo+!� �ȝ�vdm���>rfKY*[,9&W UZ
<%�~E��N��G+7�y�Q�qƮj����{YC�F�ɔ����}�p���Sn���O��U�p�<Ϋ�?���IB t�/؅��]]tU���l�|�Y؍`��'z8�l�9��*iHz��| �8��Cf��ZH1����gWь�7D��߿���|aaa�-\�>�Q(%5>�j���~Áv ���,� �q,;�1�:����=�z0{lcgו������(�<�bQ�}>n�Wh����NOg����6�D��*������9;ϭ?v��^����}$��L�D��=1ߟ�]r�����qj�+]��75Y����߀��-�Q���۾~毞s��S�1���0�J, �3ӣV��I milū:�o-�5��0��v :��3�2�K��u��_�������]W���Bi�z��/onn�lR�D/��
�L��Ngj�?8����ӊ'0���֯?���6dD��9��.��evD�t<������2c\���^N�u������_�Vd�������gZ:w�,7ch�M}��� 3�'�z�B�K��o��tqj�c�N�Ne"b⡄g2�ܑ4����^�����4#���k�u�v�O˥�O�+-��v4��;�Z��'��n+��K�(��_ރ�ŗ���ҷ�����R9�GY�B���`��D���GP���TEt�����e����l�+��@a���*���.uS��^�R٨t��3������|L�:m�9"�o�t�;���>w�V�������	d����sAT)�������_�x`��XF�R��,�F7^��7�+��0�Ҷ+��>x]����$v_)�U�(�Z{/*ޅ�LHF�oe0r�}�VO��L��H��m>��R�'�F��}��-�j:��~%=$S�F[�F���T_�Ɍu~���� V4꥓X������L�E�Q��:�Ζ�ɼ�KP�t]��M	O.`�999A�*�48CV$='%��C$��߿�Js�h�`� �R�R�C�V�S��LŏF|������N%<`����� ]6ֈ#KV22���u5�+7h���G�4�¬4�������ˋ��.&��Ђ騟��.3­�J[r��"R���z��B�����J����M�	=�o잝�D�\C�*
(e���^ԍ� �7X~J�Y��ELLNfl�����"��Á�4;Y6in�F�) r�qV�zV�m����_���j�1Rb0�N3AW�D�;@ݡ��_��~���+o|Ž�v~,	���js���|�W������'���Gd�ם#�,N�5~��"���<ɏ�����C>2��������A}}j����I��,:Ҽ9�����Ze@[&}8��kv�H��$�WfWx2�~�@K�u�m�|�.ي��@�:������04*�w<�k9?���Γ#�g�g��� 93Q��E6r 	��|�Ao22���]#~�RD��	gs����oy����p[_���<�w(�M��Z*Eܧڼnﺳ�HL�Y[q�9�/�M.����Q�^�,���E�&ƭ9(&&&�(�zEr�A�3w6w#��͍{������ R�����X��(l^E����o5��	���x�v����(dmw�d[�Z�6C��Q�׬���F^[_��1^}O�;����m��&VP�?�|g�[�{��$�q�P� *�֟�yFf������4���̌ #����������#Y�
������Fݗ�4"���}�M��o0���S&����Y�V�＆ګ�6t�����FD�c@�-j�kgg7]�*����+j����/io^�nʡ8�J0�1���m�������*k�ֽ
�L�����^؃�k�b�^,�B��ONҼb�e`���U����	����(���Eˏ]�����o(�F��7�H��+OS$��I��|T��ֈ���۩3K��Z�����I��X/i}+V�"����J����c�<��{��ؼ����>�ɨ�yYl-��m�Tu�?I.Ds�#�y���H�6E>u�� ���	Μ����D@�xCCC�jZ�sN�H���^�ϫF��M&Q(�YMMM�3źY�VHjQ��qx�[?���w?��T S�B��e��?;n!i��g����|���ů{�v�A��&S�j	�R��/Eg�����!ׂ{�h{))���mC�ߥ"�޹Q�f����0�%�CU����*�!���?�����E�0��45|�3��IJs$�l��s]��b�C��ÅI�Q5�[��?4�8�p�nE ��_�W�!)Vn�@Q�z��Ow�<&A����h.���ܕ��	�u@D�$�;�l�b�/?��g-��,7���S0W�>�� Q��=gK�p5Y��Б�������oj�v�WJJtnO�\cR��n�� �թC�e���t\N�_jܨ�����Βh?���:ktۀ���d3"�(����l�+�	�Ό����'�3mx��o��TJ�y�",�o H���1+��N)p��
}W(�Z(]��ېВ����0��@|���n3h�e���=*�1�O-̴�ٵ�ˠ��z
�I$T���zRd��RP�cz:�
�r�F�0�@9���?�漊�~R��PVk�K>��Ao�r�w�P/@�'�I�Lʳf�$��v�'c��дi!�y�(��Y˔�6V@-��ƮF����-�ٓ�T�>�^ QS�.���zYN�888��a ������yآk�ǫ��Z	f�	%m�ī�PDP�jJP7V�'��c��J��0��{?����v�o����j�r�I�4jϓ�֭[�jP"�2B���H���[�P���고�W��}#
�+���gw�~_�C�8�%��hvn.Hx��ԝ�9�?�i��}-~pn]U�����X �{xH�O�ɘ�S��e�|��Ņ����d�A���Ž�m����-��(-�Z���6��^�¼����#sf���D��O�ـ�K~ͫ��'�0�tE�b�V�p�a�,�ZKb(وn��C	����b(
��߀�X�b>��M.���Elsss,�)U~*��xM�)�W��Ӄ��U�<�AO�q�Ƌ�B��=���z��H~��/:��T��2�X)o�ÒJڲ�s�w��Q��>;�็�*����$x�n��^%A��]�g�J�� ��I=��{WKMǢ�rƾ�4�Xj~X�JE��?88�z�S\O��S�ea1�P>��=����=݆�)ѥ����!�	�&�\2ׯ��.��Ȃ��Z*��_F_l����R�^�Vrw��T�x��P:Q�(��ׯ?�ǖ'ÅN.������t��j��HSSs�3�֮w����v1y�2�:���QkN�^5 �z�,�^{G1p���:�	�s��p�V�z��}��f���Jj ����x�����0��/ۍ����S&�[���cK�Ov=e&x����v)7,�%�?2�\�Zf�'�g��Ҕan�|��l�����8E��#v����ͱ�n��4�r����p�J��e�R�+�,%$2L�����]�a��b�t�D�� �{s
+=[^(��7/E�Fq��&�̮&@�զ̈́�Fz��PW7/����\ V���?�1D��J�9XYAg�����KO��fB�>�T��]ξiK�0��"<��������=;>6p3��|/�G�P�Ku6Sf{f���&=�~d\K�ƙ�0���E�(����E�k�?ᛜ��+�����;G��`�U����N�5~_P�Z�m���}==��ʾ��RS[{)F|���<Wb;�AN�v�YW�m��kW+�X�?�,�k�Hz�H}5!$�������f��ܕ%ᶢ����F���[P>�oM�+�Ʋ�Ȕ*�jd�8��<������j�fĠ{!�/.v.� n#[�a^��&�/���)�	�H{{;z�5荬�!��o�udۧ�� ѢW���7�⋓oƿ�����/GG-�-f�ر�,2�[�d,���$X�D�Oˮ+�)sz�fr`��m�w�u�l���1>C������"�H��z7P`�ﶻԧ�]�
�����9F��z��l����lJj�b��&������(o����Xu�?�l�N��r�~��LNZn��'��Q)<~���%�CM'��C`'����=3?~Tu؁�;��q�,�od� �xE[��m�^��?'y��@
Gp��8j�U*�!�Cl�k`1����sqT砘�t��9:��/�imc�#]�В:&.��۱i��2L��**��B���+���&�P\��fc ���5z�y#�����4�ty�ْ̆�g�PG����_}�k[[uvx--�Pi����>h	�/_�_�PM���=7'����G߲ZEe,)ѳb���y@�3��I
d�Uv����%��v�{oB5��<���'{?7:��x��iN��&�VN��*�f�P˨�}V��N�ZT���{]b|�߿�O���1� �؞m����S�Zh,$~Vۼ��Δۇ�%A	�Sn��g��ݚfr^o�h ,���ۖ���	W"��x���J%A7�jx�g�C�)�JÅ7�_%�a�Ky�-V����1������u�.A����e������f`9h`9��D�hc�w8JD�?fg ɤ���;�ޤ�2�s��U����N�΢N��?�'`9�7�8::Nb�.�mg�v����wL���Mv")|��e3z�Z���~�,�P�Vj��}�V�ƕ����%���̧���Fi�ؠ�д6>�F��(;D��YzT����h1e�mݷ~�[Ѐ/�S&G��(~�*��m��С�-]��t�l\:I�g���5��5��q��(�k�0�ž���HT{���a����p7L��eSn����a\��GAr�S-#�v` �}e���x��϶���A�A,/��x�2*�@�e�� ����O��x[�P��8
y]�H,׺~FK6 �nhh��Ŋ]��-:zz��am~��k��^A,T�P8h�DF���L�$;f9�A\���_`��>�[X(�H�f��������<��fٗ�yu����"��tI/ � ��YHѶ��a�q�����r�4�]V��D	��N7�Ǧ�e�xY�=�u�=�5�F%8]H��k�И�5T���������T��˩V�Ԙ	��7���G�H��̒r�9;;�<�-��8�d����#���t��A��%�%fjC�'VbZ��Pzz+�������xq��5��u�@}{Ɍ�����l�bL��;Z�ߴl��.k[���9�~���Ǟ�����ӧOWs �Q~[3�Cȶ��ҵ߿��2KIKC(v�6\�y?����/�8z��
�Y�����YPD���$�(yK#���;�~q�s�� �o�L�~� ��&�At��t��p�;��� ��EE����@�Kژ��5V�A�2�� ���^�,:�se���Γ���X��>\��@˛�!7������ff�r�qTF��@�e�q���&:�y�?ll�����ŏs�8ɮ�<���4ǫ�@	��I�+]�2ï�	YQ��QMPf�vi�s*���wParQ�D�6���������/����8_��y���HLO���F��^��E���^��~^��T^-���8 �|?�����l2v��)�d����=.�#%2����N�7��V���^(]����`%-xm����X��( �K	���u�Le�(�9]F-o�d��o�R�}ʀ�i��$����:�n����u�P zKKS,�i	x����nz��^���lO�Y�A%VtιT�X�Td�Q X6�Z�B�M��銡�U!���=)Tǫ�|%��<v ֋�s7h�W�e.�E������v����딍�e�^5�\F3����
3?��j�w=//��=7YD58��Ă�� �y�w�t�J?).�.?cz�t�z"���6�iK�\-�~�&W�",I�F��g+�dn�������<R��7붦����Z�bP4bK/����m��_���%�d{.�j�������[��w�,��@�c~�ը�-��B֧$a�c��C/N�f\��j2�h�\��?�[�t�2Z���n~! ��m>p�$�*a�����6Ƴí�yk3:@���ϕ�˲���9��ΖJ�w�����=�
t�����|��C�!�.�}��g��U)T��^u,���P�𫥈�ee��ۉ��=e��f#������^���bĢF1绯�a|=�������C�� Y�B����~||�d!�>sm�tj?��% 4p�׽�]\�q�B�&�Q�L��킧P�)e�2Y��U�mm04���+"��l�VY�)�h\��_W����I|��ʺ�>!��ߛ��o=��+��PE�����`Ȃ��?����r���EV]]��r��o��V��Ž�|�\�_�BD��*����ޚJ�{�O������J"�z�򴼝Y@�@{c$NE-��UX*�Ѓ �;f�8��d~
����"9�'�Reɯ<n|6$Ȍ�N߶������1�̤���!ψ�������)j_�-�?�-�l�H��UM��ppp$|��^� 0��9G�xGa�ez���#���DD�u3�(��,*����ؐ�;uE���*Y�;�/N�I�ڋ�<��w/|8�*���g�����X��(�a�3��lv喖~,+�*�1B�o�$�:C,yq��[CP6��P�F������|�����ՙ.��/"H��l�m0AEto�_R��}x���U2ݼ�ȧUB�h��㳥�x�CP*$ZBYxV	�x��2�>��p�ja�`y�_���&�o3�	���9sq`'�'@)��9"��)������{��L��V�:�m�٬}IO�%��7�AYf_�mď�3��x���H�*[/dZ�8$3*+�����N� �T���{���-�n�/A����/n��\I��F7f�xv"x�ԛ�W���P�Cz<;�v��ni�f;�Q$-����I���f5��(fvv�;8-)��"G:{��tM�c�1<v(���痏.i��!3[EB��/\Mz�l;���ۢ�6���/��ý8���Z�v�E�Z����ۡq㮌e��N��r�-���FFQ�1�pN*��|�xUJNF< ��8��(T{�W.t�u�����
���%��,�g�tM3W׉�3���4����N��fW��&@��yHC���¨�WǢ��[ﶢ������ ���#M)<��@�5a�.~,!灑���}W����N�v�P-�
N�*.�g�w#����8����r�y�^���#��oWȑ�7zZ}8�?��n<;^xў:���Xؕ�!(�k�;��V>�0�Q+J(c�iX��}qq��qy�D��,`sG�ĭ$���*�SI� |wf��0y���i9ZZ��[g����u������ytK�p�` �Wk����"����<ɀ:>42���[~���<{�z�/�3�h��d�wy�tEؼ�����c�KKźD�&�￵7���}I.��\1��א�$\����z�5�[���}I�m����2�����ۊ��A�ug�6���� � 1Wz]�Wײ3ԗ�x$L.��^�%8�h�3���i ��XB:@W����bbb/;���ԩ6Itu�=��Xi�w��g4_�M��y��#�������~d�n������cI_�������}���IX�m�~e(� t���{���Ts�aZ���8���		t>��^3��#Sww�������0 UJ-�!�}��׍�ЅE�a斍���M�,��WG}H�!տ��h1�W�o��m��s�M�2�I�߱8�ߩF�s��J�����i��P�,y�o���8XP��d�!�8��q@�h�c�˽�q��-r	g����Y���9�0����=Y�o�u�QBSài�ܚ�Q�Ȅv�z��{�+�:�h+��	F�\c�/� ����#^)3���P�/�y�Ih|��kG�moo���}������f&��~�����sP.���e\�_���ի0����׽��خn��J%��KO�K_8%cLmneYYG���`��* :O�:[py������n�A�
R��;�>?.�=�-;iǦٵ���H��ܔ	�P,�g�����~z�z�vC����Prz��Ol2Ū1�� �,N V��)�j��+��A��޾J蝱o"�c9�����A65�5��)��;455����Fc��&�s���C�{��S�w,��aWN��єۂM �y_�y�E�M�gL[CZ�O�5�8����މ���]��@�]Hs�m7��]TF��x�9z~z ��:>����J��6o_��E��2I��z��#��Sy�ұ�&��������)	%�ܛ�T�l����PTѹ�mX��R	"R�_����V6�M���	e� ��(/�T���7�/�%�'�po���h���d�I	Xk��L� �'K&�r�s��6Ubf���.9��������>�m��\�����`oMtWuAQQ��!�~2��?�잻�x{c�����d���0��Ҳ��� ��Wj�V���g̹ڌ�]�Q#��2k�*=�Zu��VVV�Mmd�zhh>���v�� ;&'�����8�t��r����u?&��7ocI%��������+��xo�ώ
лi�g�7q�g�ɓ�B��i�	�`���bg"#o������X��O��gQ�V>����Ο|������VTV6��^p+ V�^��@�ul�o�Xy���� CB�#3 W�w�B4u���Z���q4�p��$�A/:��� �0�o���� ~��5W~c~���<P��Nfv�&U�ׯa�&S�9.�J����YVl���=h[ށ�S3�Kx��ȓ)A5E�3�SzQS;�ؖ�W��$&u/�C�����@�w#���&��$a+������{�cV\J2�l
���[B	�5y��|0ixI��i���U�n(��TÃ�&��n��V�E@4��8�v�[��lH��v����x���η2BŜ-��'&'S|���锕��KI=��P���`��C8���M��8�{4,
�2�]~�+V&���l�s����~s��wש��|K%�k�C�)�����F�QހX�ʊ%��e>���E���$�R:�뿺���_�8���t�"�Q�� 짨�a����?e��r*
�GP�0��v񭌢��������D�F�!�rP}h� z�za�!�$���!Q��f7o"P0�6���n�ʕ�2.�f�q&�T/�7*ۘv|�Ϫ^/u~�v��ӻ��Po�z$}�6x4�%�µ��}K��� ����U�vB��&.|�WWee	�یC�ǹBn�m��7r��Z�݈��ԪPƧ�M��R�C�Ļ�Hn,����o���+������2y�������0hr��&���������������y�FZ������U�XLB�%�QR��EbiiY%\���%TD@$�F�A��o���|�=���>3w\�u��3ϯ�ms������ș7$�����6m�أ���_���8�e!��[�(\R����� 8;:���?���j7˙�|�'_�xhc��;\��i�;5� ��Gך��6eK�C����Ӵ����l��!�2�>�u��_`g��{:�T�.��#݉T��?+���UK�y1F�����9�j��6��̸ W�^�pƦ(Z��NI�X���!?�"Qb>�su}u}��kM���k��,���=���9
����7�L�ݽS$x���� �J33�u�s7��(�QX;�fP�7�ػn�'�_��`�	�\��E�.y7,?��t��5����(���=��!/�nh�:���V+.>#����m`5�3Rܳ	^K���]�9R�bee-q�V�nTϼ������{*.���}��3��"�WpL�bV ��q�F$
�5�iBd�u���"��/���ꆾ��v	_kQ���Oo'>D�y��9�X�/bFG�&��)=N���~�����u�-�͵�Q�hN�c-�U/bŠ8����[7���⎦)�qQ�_�C"�4<0ħ�8�����[����_���KƟu�6���e���d��(�����nPC{��� fq}=���/�{L�����j��&�C+����0��D�h���X`�rU[�;%K��~�Y��G�mx3׶G�~`��Q9Q<Vg-w��$���&H��u:u��h�5 &é���+�ۍc��kl�Y4G�"Q��G����)!P7���F'��ӝ��������'I�b�@E�"�d���}敢s52=L���W����mEM�*}t������c�rB�7C+��?�؏�!��}}}�G�����D�ء~(M�w���gE-�@�ytbNEdq�s+���K������nN\�o�t����4��B�}�F����w{�g(�
�{�G=3*����xM���C�]�����W*ؔ�ۜ3�#���N�O��8��&[f�d��8�6w��^Uh��~yy�9,���ף,�lS�;��/�� V6�9��n�F_@�]W���9Ei��8��4��H�����WA�� ""�U�`��F�h;T3tݐ[��}Z����\��ƞ�'u���<��۷ob
��S�Ȟ��ܥ��u���j���*�ٔ�3����ܴK�d�V�	���Z��*�Q����`�`	"�|pU���?�:WV&0��2ΐ��^H:9��wlQby˳Ĭ�P��9g��]'���B���AkJ��b���ۉ�U�B��dO�cN�[ݻYu��ne�?ee]����t-j��ښ����ʟk��1���+���DrU6�`|ϴ�oy�(9���%FYQ]s0��瞴}�[�egO̬K��Q]�L��:����:�A�5[�=S�uޛ�+��5���k_�/�@�0���L-���X�Q��*�e��5s��ӭ����qݯ�|�o<ײ�}����(
��;e�f��VIlU�9�\E%l�Ut�l���c������px��ghH�A�#��?�M|+�#.��7�JWُ۬�qh��^����uզ=���f��m��bɃA>��7x��S��kɪnI�xv��/?O�9��Et�_@�4��YZ�u}���-2�Ň�=I�`F=6MῙ���OW 5��$�BD���@�h,t�אD��L�Ũ�)Ĕ;Y��.��rĕ���
F��=s��^ �����p����ѽ��_˽i%�H�u�2b��q�
�p���뤼�����1�rm��|��їDj���3��y*�5|]�vʽ�J����c�p���������$%NT�NO|zk�B1���\�����&.9��1��B��������)����I/�>��|x�;��)��}���Yh��CKP��Qg������Z���(h���$��٧v�$<�l �L�V���?+L�K���!W�a{*xe��|&�x`Q�\G
]-n�_5�X�IRe�>�ȕ!\�#�]��D��弟���:he��Iб9�Pkjv�-�'���GY-���:3��͕�Ks.FN�l�������(�Я�����	���Qbr�!�ژu�,V�NSUL�Zd/2�+y5$�:R�[���۳���I?f/��*Z�S��^NɁ�� �`2�{������	���>S���+��#�g�m�B����7�����O��h�/Xf��6q�I�#Df�i0k�^xz2�YU�����͛h�8��d�����y�����sO8/4�\�E͋��#�/�qN�ErY���G���rR(�b5��Q@n�������u>d��䆎Rtww���u[�z���9�c�l7�wzzV�]y���JJD`�ij��R���r.D�����a娰�� ��E��O�k����P�k@�vjy
�ze��z!���x/�]���uDD�C���a�AP��`����߿o�?�R扽�M+�����:�Z\L,�SFn�Ewn����˕���Cfw.�:�T��X�UG�j����L6�S���I���w�u
X�~4��^b��/�93�/j|�:g��_~��1(�f��{��U�
��>ܴ�����C�D�.qƐ�]�N;��`�Vf`�d�����~J�Vp����d��h^�[�fv�{s�8�W�0N��ۄC��b&��p(��0���L�}���U�#���Ћn5��G��0_�}�a�[���M�^8wJ=�ڼ'_�-\�?�&-]�W׮��ၼ�=u_��9V�.4������6:u���d�W�ݧ%.x^I��hת��>��يk�U�\����U.Wk��~u�m'�7�7~��h�0<�D����P��h�q2('/��T����%N�����c����S=���v[������y��K�r}p�g{~�M2(��☧�N1Wfxa'���2��.Au��s�Rf�Q�e�=BCGG"X�*FD8`�ܒ��P
�.%��~�_�Xk�}�U8Sc.=��j����6on:��}d�&���[�9�~vJ��[�VH�����P�7��t׌{ص��Z�M��l>e
٪|��Bg��;�T�M�G��zHc�L�Q��خ����C��G{�YJ��'��)��
����;�f�G�������?���on����^�z1��Z��G��cub>O~�����r[}�!�$s���6
~n.�n刭#�HE�1M��ٚz�bs��EӖ�W ��M�����/�G���)���be[����0+^����Z�!�B�%���s��Wv����b��/_�����<I[cw��Ů�	�Ŭ��X�Й��A�;�7Xi\;OC=�8��򞟏��x*���=�[�o�;��Xr5��(5�!����΁�._����VW)�A?�j�'�ק�	S4[���%��;�%-}ֽ�)#9y�qP�Ҵ?G�k�.|��;O�������1�)ֵE�>}z1V'.��Ό�Έ~������2�Z /6�l��������dx��e֡���_�u?5@6�+]���HA��w�?�jc3�d�RnV��,`��M�8\W�<�L K��L���^���S�W)���t���@|��I��x��8�ӿ��>S���Bfouy0�|�iC��kZ��ţ�����,�w���w�\S}�b��?.s�?��UIz�c͇LL�	3C�^����-���pn�ta�ќ���P舃�߱$t�b��������h����������g;�t�^~W��z>�.�@��~d��3c�C��VGj�{Nf$��<)�z�nϕA�=mo%�O�Ha9�d�^V�N��G�8^ȒX�/��7,~���$&^����N��1@��ǻ`x�,,�K�}��$P�ȎcȞ��+#)�|�pu(����ג��B��}cc���?���7��w�6��)?XCh��ϳx��:�}w�j4��p2��C=+<�ַ��Jr���L;cA\��J?�Njp����@�Yi7�}:9q��DtF���[���'�ok�IW�%}}���Q�����rP����ōg_ X:-���q����b��Ђ�G|�&|2dd�TX��1Vɵ'��<,; Nm�Ψ�}���DI��觚����QgϽ��5�����z����@;���H��0t
���ts||�V��� ��"�UE4����}���'�R�y�)����������ټ�w5���������/1�r������.= z$ ��f�Q�B0���k
���<9PM�4��J��鄙�ڭ�����od��YV��9��J F�(��U����R�?��LV�Y�B첨�O��o��C�7o���QRS����}��]����*���⸐R��K��ED`p��F0�7\�T9�Kf�L�#�|���_zY쎹;������N����Ԫ���k�E�{��1��uΠ�?�b~�����gD��ǫǇ9�r~�![�vUU�;Ȓ��/�̤e#׷|���, �;x���ć ��	�q�0mL',���%�pyej:��	���KH@|�ƍ@���ﲈt��rN��}ХuĄ��y��[�IZ���R�ҝ8��v���/<hrKO}��#'>D�E[a�[Xߚ���R?���1��{37��o��H��]�{a�IIL����B����5����k	�`���2��R��B�8�3��M���Ukɕu˓�ϊ�Y�[�ܑd�'��0�P�;ZB�>rƔ��_����4@��l��,x|5e�\t��v��@ �������9��ee7c�Cל�׉p�%�B[.�7mɀ�}��ة�rRn����g|O����W��5t2W���7��|f������l ��<M�]�s�������k�#�~n�����z�C���y���GT�o��l��QP���nCC�Y��d۶5	�+Ýdq���>�E����|<�X�j���x,�[J6g�Ώ�^.�M��}�� �t�C_����@;2���((��M�#���J::L�-&z�u�)���xQ����:qEX��9F�,�q~�2 DS����g�	㐗��>����Vn+��zǑ+9�8�6@���WD!�c0[t����-%�{u%��J�dty9=��1y�~���Ͱ}�s�x��-S_�AQ�
����M%�����P&����b�;�V�'fZɊ�ì�;~Eo�)d?�����	oʝ@n���z"���卉���a�	"��Q���������&�gu@�<D''��VVj�~���t2�B��=,��� :�jv��n�hI�X9^�}�Z����!�{	M�W��l����g�xxH�^��P��B	!h4C��l�o��L��[��V�G-� ���U�'wLǚDM\���ؠJ��Kʴ��\ f�����4
�0ď6�N�C�ʓ"O�Aؠ��ո�T	t2�#:-d�`8���R��{��"I�Sp_�f̤�Y��ddv���"?��[������_/�|�B_�m�����'w��)J��P9d�����s��>Nkl{K�.)��u��@�a� ��F���T	CQ%%�_��v�)��k;66��8�D!�k��9�H��T����D�"��2���4��z�0���*��[�LeJ�����5�a��8)f��.K�Y{KfR���|�<2�1�u�s��n�/��Q���HD�H�B�3HeE��5]��?�?�O�9y��[�WOկ���VM���v��S�7�O�Iٙ�99:�6 �w	F�R�`�34�]rMl(.Z!'}]�)�|�� Q	��j�rs�|}}�Y����J�gP�F�f˥T��z�����[N#�J��'lg;R�K�dxx�!�Y���� HT�`c ��Aѭ�������^���H���(���f���eu�â�PTW�)�[��eܰ}�����Sr,`ET�te8�z於��4LU�Q
<q+�L���D���`���L��au��io�%�eDy��E���y �i�~�K�Y��z��e����x3����픣�S2e�������NM��{�%˝�p�c]��&�r��5��R'�>g��U{g˪l�O��{�7���۴+a7�{.�W�������� 3x���g-|*hbe�?�B�w}�ˮ2�*F�VZr�զ��KC8)�������vkOZ� 	�?��5�����OB��40�Yu��/ڭP,�����$�n��βc���'O�
���g��l/�̝�P�
���ǻ�
��q�0�=����<722�;�+�h?��E��iB�G{鋗�e�aݔ��&�em�ƹ�6<qR����������W�X�Е�1rB�{�-�7� 1���t��8�+��@��Q ����sE��t�픜+��1G�snK��un=0��B�� �%�����%�+mV����}�g?+��i=��)˛k��GZX��u�w�|�{R��D�z +7�qT��U`�PZ�r�����5��#�]��#9���-יK�d�g���?�1�
�'��2�U��j�iw7�E�3� �q�S$Vlj��.34oP�kY���Q 蹱�6�J�Ó���@�ؑ����ޥM�/��K��޿.<5s�rC�D�B�S
y���1Q��y��Vw��޳<P�%���� �Xna���E�bKR �?f��Q�9E$�qVnn(�0����4(Ea[� �0gn��K@]b�Xz��� �9!����,ȑ4L�ZI��.���ك�8�d�ȿ#��:s��~�t��6�������>YR�y���b�)�L��"+�Pl��h��e{q��7�M��n�jq9��B�:W�Ԟ:͈!���Md:ʢRy-�l7���$��*/兿�W�-�JK>,G�g�9��@�	�Z15ܬ�C!Fx�y\��\�ס9�;�ͩC�*Hw�my��J�^
	3M���j�9�i�=��>��u:_�m�u�c�3�LwJa:�qc�$�/���8��n&�Kw15�7%����X�-Cn������(# ߚk/6wt�g	R��$�[�W�L�;�/���g_W�lM�S΄-`��x0��?@��t���jz�g��nV_t�d򦾯o����Pډ�&w�J��jxg>�~;�8
��طL>�k�
ONN���}�hh��K�ZxeQ���w�-B�by�.��q��.6�J6>�(MW|�W�&��l/_�sm7DD�.;uO��)ٵWb��|x��C`�A��7ZP��6�05���|�	���K:Oӈ탫~+3`,�E��Nۍ����T׶Վs?ml\=���~�D6*)�Bل�48u�����Pc	�2qf�κs�fO��m�-޹��tȓ�ղ�����zeX8��B[I�IP�ɟ���q���Q�<�v���$��6Gjׅ�<�Ɓ�l9�vRL�ƥ�dO�(��_���j�����W.��U7xѣ-:�<)��j�\GGu��N&�h������oC處�Z�A��}�<�͑$���Y�>W|{yi�������>�L[Z����S*�*�J����k��X�V5sq'����J��� F�
$�<q��Ԡw���Y�-V��Ds��!9�����#�C��!z8�x�w}jN�����z��(�<��fVV䠐1VJz;Ÿ��!����?nbJ��5I�bo�|ݷb�@hCi,{kTS������M�D�2�f7ݫ��>I�F�$�e��w�j�y��
-�2���_4Q��oh(PP4p7XC.<���nEb
j�U��#ث��7��ˇw \Y<c']��ʻ���9��B�کo+{ͬ:���Է�A�fu��<�'�a��zEy��YKF��.4MҨ�cj�8�v%���><<|�2�J��ޕYh!������f�N���!+��0��Ŷ�I�)i�Y�]ر���y_�(�)���|`F�u��Lw�z��V�ꍼ�,�dn�HF ������S��
�%��	F� �6��@�� ����/(�҄f�E]�a��E�)�����`��-�0��$�2A�Q�A���u0&�B0���X�|�m�@G��_�o2�{���J����4F-�|f6���{(��k�tL �������̔���M�_�pjWЫ~|�}3,-�]	aqc���?=g�$��=*��_�_}��/2F/\FO~�P�H�m��9ֶqTyW������ì���ue��b8t���ڞ5�h�3y(�CZ�X$�;�@S�ҵ�����>D�������$Rְm2�u k�ܡ�߉X۟����rk�g��+e��:�{���(��+<)�+Y?�Ƿ�zG�"��H����,�R7M: v��wi�d�i��O�v��Vx��l�����ſ-t:��R ���3az뎦k��^s�������_
8���}2��;��!����
U*��=���$A��]�a��5l��T���W�|~_K�`8#�`.�����E���@�z&��������C^!��Ti��]K��,h��C�.!멠������I.�(��@y��@�
���5%���=��(���ږ�S6���=�ޒwxL�02�/:�JQe�tNd ��aԡ���r~Չr�	���.�º/ ��<:a�Q 9��^w��v�n\	�j\��Ȭ�N깻�g�x'w+%zh��-���G)-L�̨
���ٮ�2�[��D�#�G������G��.s
f���;__�3��U���:A�Mv���U�5
)��PW�1+�E�+kL�L��e	���h�Ccg����f�Q��~�ÿ�;�b�]R�Md���J[fVL4;^2,k<�2b$��)]q�5��黬�ǌ����+���䄼�����b��3�� �'u1E�B{Ԟ(`T7U�����xïL2]�S�3�C:%�ٚ�����'3�1��#�S]�O|��{�.c��S!X��q�Kz����-��9��$*�	���E�ՠ�YU�S�r�Y@�Z����k���㈑H�T���V�x�IW�J����2�(q�^?<kJIM����_c�L����s���.�Fa?�orR~���$��Լ��ҐH�kΩ�b�������0��E��}�����F	�Ǜ����.��ﮧ9z��
�q�����q ���1a���L��=<:���{3=mJ���'�B�� }WWWnfJ�SA-�~���� ��ǝ��aHhW�f�� ܿ^�����U=;��ïŬ :��L� 5d["�j����J����,��+��ke��¾ifъ�*=gL�z\�%���f1{6���)���}����-#�����@X0��}�{��i>�L�~u���. ���Ӌ�ט�i��;�F�^�w/N����>��\���@�q.��G���'	��u���v���.Rw|75*h�K���-���#��E��(���
�`��� qwP��,�pk"��T`�P��2Ӆ!���d�����$JOO������^��ا~s��5鑁��\,m��������F2޶��w�tۼ
��fYy�	�zI����o������=Cex0`׻@���m����"S�VT�~�B� TS�?�C�x�5tt��Q��G���>�(	R/��^	E�_?=�I�/ܡa�vط�b!�\n�+��B�'%
�����߷�0�}3x�� �[�@M�"˓��6�>���߮jl� ��Cr3�`0 |M�����p^�0�}�pe�}5�? �ta&@�g=%_r������
�^���.����C�	��M��~��{���.5�i���ف,s�K�5u��Yj>}�_ ��3a�v�2��-&�1�2{dx!������qZ~{d�K�g	yc �#Gc8��W����hn�bQ	���c��}�K��"��W:^���G�m��K�73��2U���9Q2���~�Kf߰�Z;	CY�B�u��K��5���UxݠH>Vԝ��KX����L�~(T5��xF���wH0k�Q�ŌJ�Q�,�k3��י�,��}I��Q�a����JL��X+�W�q�UKWS�BL���ߙ�
�������a�	�]J��yэ��y��DD���mn����e5\���_��1&|�E/	{����ѝ6ɐ�o�wHQ�.����;�[ �c�k�ߖ';���*!�� �J�YYW�߶\�8B�����(���7���ַ�=�ըޡ;	"k:n㳲s��_]8�?I��ngptP�}P�F˛�*Љ�m����8U7'��'�B�|&W+�'tpP[�*z�%QJ�B?�9D��M�`8���� �?{*ϓ�[�w^t�������q���O�j)�lIB�>���S�t��9R]X�[�%;�ῢ�;��PhC����JL�w��4��W����R���%=����P����\G�`�$�$w�M�~D��<�M���'�E˵Ԡ�t^��b��=Ά�Gɉ1r���^���{t[6 ��tr��?�&o�ὖ����'�(%�6�n?p�\[���/M��u�A���Гx(���	�ɔe�洮?��b�Cݑ��ۃ7�2c��l"ß"�~<�EpF>	P�uZL��0�:e�Hq�T��3:��t9�Jj���K	��}���iW)��g(�H�ō��kz��A��	��o7,����O8�����"j�Ēl0H�=����T?}��u��i����|+;_3OS��q�Q�wp�cY�j�L
��H��\f��L=��i��^!���!�؇ܩ�j@��ߙ��ѣ�H�HL�D�����~�,j��+�̕�L�6*�	K��<�B�f���݀����UYe�fB�i0��w�H`���m��U��W��d|�2���}����x��<��KryƓ�B�m@� �NV!�-R���@hA;��5���0� �����՝_�`&|����������Z�7٦%F��b�Ն�����]�U͓�+�B������$�Iﳍ�ʳ�'2���MWCN?����%�����ZG��Ab�(�9�j#%H�~(�����'��z&�>qUz�}V���$�z�o��Rp}��X������:���F�$ӷ=O	 �����g�UW7D��	b�w�Qwޖkiw~��	�g1h}o[0Jn}6��eA���(�\K�m,>>�˲���0B>r\���K`���X�z���u۽�a�0�d��p��5�tq���Ė;�f�!����~���]��B7�$��Е�&���_0�"������?�r�k7"�mG.
�^�8�����y��
%(����B�=fh7���l���Ͻ�z����(F
F�[*q�O��*(Eo����~I����<�&i�؂d�3��:�-V=��+@��Ͼ<�>�� c���9�T��³���]&��M�@�"��	�pQ����ix��uĥ-���)���C��u�+E��^���Q�ڵ��B=_l���(�Wg���$S/��S< 5�#�ߖ���L$�G<��,�?hu�%m@$�?j>�!o�SA���@ ��[[葼w�Z�
��JL�ԛ���pk��?���ԃ&����_��\:uc���% ���#e��j�������y��q�H�U��ғI?�p��L'��{|)��	�EsT��V�ћ��}�	]s���K�u���n�b�&�X6j���k1����w}7����}��Cd՞|/���5�A����6&���mL�\WvvkXN6 ��h�
@#���N��1���W�f�Z�~���;KvՀȊ$�^7k
L@�d�2/./��3˰&��\��5c�?n�4*g,c�|�ˇX˂�����A���4qPOS%�P.W��<�#Q#h�������נLF�:���w�u�K�y�/�
-O��� ��1����De��r9����r]��`� �	�(f�����Z<	L�aYǌ��`bB�����ެ��;���dtĴӨ�yv~
�w0CL�Đ{�zq��qa����z��7E;%!���u�nz��|5.
�|�gf�R0!Epk�,�C���|r�/&u�OE�)��މ W�(�;�W_��}�<�'x��Qdh�������l�s(j<��4=z���$����h��9���z�3}q^>�7^�mLr�4�QG�f�A��kNڵ"�p�Ԥ��Q�0�u��`�,�f����C7A�1���Bnڋ?^�?>y0|��a���k	�����ٽCCd.qr˵�f.I�z�1�o%���3+�^��!��M�˃�����fz�B���ȳ���ǿ��j�(~�zE��O���tp���(��Fm���K������p�?e I���\r-����>�7m�巀�{�|�x����UW�V[�^�VL]+�����b���M���{�14����c:�����R�1���j�u�ݜp��:�$#p\
'�������mr�=�X7^���#�	�>�h����m�B��cqKru��\���-ï��� ��+�aQ@����v�Y����<�m���6;)��-/]=�\0<�� '�(�#�RX,݀����`:^a_QQ�kJ��=/0��h^`�5Δ���F>�g�#m�/<M��-������ap�:v-a���o�x;�$���~��%<�����G՗r>�Ŝ>;�.N����	�3�c���3��P9�D<h:T`@h��*{�2�H�q'��MW�Y�)�t�%T��r���@ݱ�����hDh��-� 7Pāh$w��a0�I��Ӧ�fR�A[�qu������������E&��3W9�ʫ���T�X�4�e������n)@ \.����oG��K��c��I#Q��1AIɯ慪�)mV�m6����e&��%�	'�5��<��~�i=Z0����h�,�@�#�P�1��.Hg\E��ች����w�p�A���Qa��?LU���Q�f˙�K�֌@`��b?��._o�v�J_s=��3A@0��#�?��z��q�����\�az��{r���-+�F�/`�N?�&���}�ۙT0�
�T7Za��V(���R~���֩����u(��J���S�8N��_IN�����dj$���vg�qG4����ZLǤ�k����2�~�W)B������9�AeF�aG��.�8l��E9gɒ��L$I��b!��Ol̬�ph���F��^���S��Q��n��S����6�Hî8�b�)���7y*T�$d��7tA�@�K�u��-mv������5|�贋�'R �sw�s�/y混�ZP%W���5�n�Sȱ�������
��އ�|n�2�R`$�^�=4����%��-G튪��c
��3�3y�H��~h������'X��RY�j�oC��TG���ՐT������P����DY��)����ϟzb��~js"n�%.�\�'υ]���G(yN�{<ѝ���T���ޭ����ڒ֍����k�N�nq��:�&;�+����������*�=���(�ړ��-���9a���4r҄��͡��
�ջ ��Mwg���z[���t���M���D�y����7�'˫���%��Gۥ��d�c���ǤbT��g�a�/�p�������Z��%�p4Ù
eu���>}����m��v:���+���T���'��p�^
�vlPȋ����L�X=��T�A����ƨ�(�
�X(�U�9P�?�_���3k��_pl��-l ����$� �'�*�d�������â�7U�n{�v������@��i.�`�8Ԇ{!q��n�AP[t��"m@�Al�ȓ�����◯����Jѳ�e͚�担.S��j�@7#1�����I�3�찚�_���k���v��&=����@��7�tknȡtm�Q9�E�W%:�Ufbi���~�ͼxc��g�R�O�Go@�u-}��}��Q�vZ���p��r�ZH�a���e�R����Sd����~N =�h����g�K�̜͆���i�����t ����=?�gģȡ�h�҅�8������;���[�����dq��3�b���9�/��=���V_�����R�+�8S�ف$sн���!�}��!.��y���寉��'�@�/˳+s�7��dF�gԫ�����zR,{�Yf�M��5 E�G!�v�{c"|�kٖ�j���z�5�=GVG���=�ח�M�իWl.5��>��T�����Jͩ�i>��Fs�u]C�')����F%V��^!kܒ kt�';�����nܽ�������6�6��c�]ϙ|��/�gg��ȍ�a�B�du��WO�9ՍC'��wP���}�,�~x'�⁏N�_&;�L��
js��y�6��N��{��3�Y�hǆ���׬'��o=�ҏV�PV�fOXx�B[�����-<�N��U��'DGꍦr��Jju�k����9�����Y(���AmŸVyac�dk�Q�/]�a�R^���e���i��l���UR9K��W�j���b����m��h��URR�K���1ͽD%'O�>���`V�����2��H����!��r�DV7�&C5�sE'���������>�IqI6�!���Z�ť|m���D���Nm�Ծ�����F�!�5}�4g��òFQ�~g	�)���Z�����52�;��r��jmUK�b_糭f��;}��mY�Y�<e�V� ������4o/�_2��W��M�J�h;�f���¤�X�:{�@�}��7	ŕ :�� ��Nb���{a;B��Н@nl\.JGO^���no��we_�����;�&���J5 }���/՝��/���d�Q�.L�={�2���4`{$����=��Sn#ME#�i�g�ĳ��!y�o�l�+��@?�ڢO�I��$T��Q [�������qݯ�#��Ɏ���^Ǖx���Ky֡�7����\9>�e�ɟ-�~��(~��SrZ�ڸ..)�R���cEA?y��!o��Ӛ��/3��Bݯ�űPo:ύj�H 4���`}w���*�OU���Ǵs慣B3/e�X�k'�x�?)e������H�h�5$:�XC��K�����SP��3
o��B=��ط�Ə��3SX�q�EY5�[1���:~���'.wr�fz;�@�Z�dBS�_��WHMA@�C���oV'~���㪺�O��.����/^/��r]�?�P��L�[dF vH 2w�� e�A��9;.%� .?+�_6;��͆ui����χ�T'''|4Z��@�޼y3�
��wU��L��;���Ԟ�WBlq�Gu[��� �Vu��+i�7'(���5?��ń��OH���Xs��o������A��4���e��a�L�?Ɍ���2&��ы��z���c烍����Q�y6�uPw����I�_-Xd��4����%5j��pT�e1P^���,c�s��ݘ�dq�� c�*��B��ҳNl��~��R�� 	O@Y��rӖ�j��X�y���;>�4MF�#*���W�2�-������>����/��t�1�$��?���D�w����a��'��}�=�w�  ��B���F��I��p)<z�DaΨ�`�L����;��S�
?'����~���� ��B�������8u� e��G'?�c�ߜ`9����£/R9�}v�;t1O�q�=��8R��]k�%/���ybr��ւ����
��>��Lh��9ᡟO׿\;�џ���ۻ�];w<����ZʐsMf�M)�6����~=���n�]�ѩ��/�9���~�*cs�M�.R��J�jN-�*\<�<������&rj��||kj���V���5�"3\~��,+ �{�w���O�{�QZ$Hg��ڲ��G�.xN�[�m�&ٙ�	���z��L�+!)���Wr�l[�֦�0X��GyP���Q��
�v��6:>���@��J$��i��7z�h�Lzxt�m!����#�����SA��2<� 2�Nh�4GT�7j^ɏ�>c�E� ��!�~�Ǻ���f�S��Õ�cu��g>���4{��)��� 媫�Rr����P��R��ʯ~"%!?�{�8E	���KSO�"<����ql���J%3j~sT��i�MA��z|��`�j&3s9vsE�(n��޸{a����[�𓒑�>N0қ�il������Z���z=P~����o��F���s����,)%�sˮ`6���۪\R"�7^��x�?��{*�����������4�)c���9�xùE��x���t�c�y�wm��=W� H�I��X?�#�*�KX����n���	���d�ʿ/�RB&&����ο^z�;  �6>,-�x��j2Q��:U�z�2c�<�B��xǇB0�q��¸�.�q��6�z)[mgP����ǫU�&���v�1�ҟ�Y�!��q�C�0���g�Mut��^H�&ʱ͹OSn�>'j1r� 
8��c;��P��zz�n@\�tx��L�5����wR�D)�yV7Χ�����AZ�ZB�¤�hT�ǀݠ���ҙ�>�d�[�.-�1J��F�z6%�S5��:<�o��5��QC~�U���?V��w>YL����|̊�M4Ǽ��uUC����%�N���|��P��z������_OGT�	��:���8�H��y	�@#Et����V��ꯤJ�iw���/_���;�#�9�C�!S�7BD�F��\km�I_0
ٹ,�Aru��p��T���[���u�B̙�2��ʋ�N�d���s����E��m�C�n�i��u�kT𣝹eұ���-��e)x�e��
�cL��&��fY�3�	<:��� @��$��F q�:��h�S�RWȗk�ϳ��j5.*$�>�o�Υ	CDU��zj���;H�a���.�W�f�@t?�؈�M]4��1,W0��^>"��%Y?i�(.�m��}-&6d�q������ћ~N58 )X^^u뎣�edh2��%����+��j;Br���� 9p��4�0^��ġ�)��Z��3>�z?�h�����Y#=��
Y�`�<&-��CG/�=��V��TV�ח�$lPkf�O���B�)DvI��I�`{�5
ݎ���/L����mm�����͉BM1����J�:J��$k�{��h1��,��	G`��+�a��/�4#n��VX���^ F�cS���m�N����n����)00wHA�֠>4���s+��O�C$�z�Qydpph����;�}�"1����d���d666�n��=�Φj�{�:桴�Ow��}���o<3�&�pjH<��6���HO�uƬ ���=%KUѭ��z��g�$�04���'�LR7���u*M>��DX\6]?�"7f7����܀�|�4w�D�e\T��>LwHw��� ))%!�tIpK���
���!��t���PC7<�����3/|�̎��u]k�u�!�m��<S�z�]A�-�#)�/L��s�2oH�P=�R+�o�6w�r[�~K��l�����B�%��-� ���L-͖���å��n����S�ܲ�Z��ÁU8�|�ӲO�%e��+��&҄u�;3�{��t|��1:�w#�Ρ��N�f�od��*h]��>�����.h�2���*��5o~�@�Z�%ޔw�%؈��`�8�k��
�q}�[��/�$���J-�B��Gr�0��]6���yoMVV�w�_� 1�m�_y�vQ�~��M&3�n%�XX~_0N�:��?{���q��6� .�=L��*��0a���c��k�{)d6w��Z�d��9�\YI�1'K���Ŗ��`_O�$���u�ę�*=l����@� 0�*r-3TUt��G{�pz1t��1QtR����c{�V6�d��*�x*��\]]}����V�����h��.�]|�ҙ��0�yM�~��e�����{��Ϡ���_i�,��
3)l�����(oun��-���L����d^�F!F��;U��
�6�;ZLe07�ǥ��.��aN��~�Hh��	����ŕ��~6궟����ӧ ��R����$uґ�ׯ_P�V�?*�����m�rͰC�~�b��M�d�:&[ܔ���$���:w�y ������n��+�T] Q�!��'܃������Άw:��gd(���!�a�.9& �?��TL���I޳���]��֙�"��!7���MϽ �&5	���=JӾel�������y\��:2ϙ?�s��w�>3XK�ű~%����`:����A�`�]�+I-���'hk=�BI�o���k�a�0@@���������l�P���}�g��Dցm��n:I��Øӵ�HRU��C��q�Q!^^�%os�<K��É$jݝ?�����i���~�X�wJJ%H'����x,��)ά�-����Ϛ`f2֨��������Jh8Q
�g��D# ��ۧ��jlZÌ2a&C�ʹjt"����b��LV�BB�rv�p��d 0`.�}H;:�V��3�x��$���,��$4�'���$i�?�i��q�O�Q�	���-�C~dU#���h�;�����z�:��6��W2습���I�n�Y7Ҽ�Њ*�@�Y�GY<���9�5�>>��\�B��Ea��ai�Z��;��_��i�X�BFmcl4.js=�����5�ɧ5rO��	�Q���iHevq��(��h��.֢䈊�+�#�:I�b^�#�#��*k�6�/�Ě
��&w ���E�� N�q�l����/��*�E���jw~!�ԥ(��Q���!{V��NDP��9��Q�D%%s�c��-a�L� i�{��a�����K&�Dվ#u��߰����^�2�S����K�� �%E��]�����#�g���߼���k����D��s�?8�ϭB@��d��v3��T�WiG�|���o����E%��*Xrw��.+㜙�y���ǋ���Ә��W�*+9>��X��:�����{g�8T�AIBR��\�V���jD��a����e����N./��aה:]B��_ꘘ��@�����o�ѹ
�����'�R�����	���9֕�io)�.�E/��G�M���%A�xP������ΛJ�S �ﺧu2[�7����|��j��$E���`V�`����^���=F�����p7b_���<���Q��y<�"$�Ǜ�j����*kE���^�,/B{05�ʴ���z_񣒮~�8r�/�� ��t�$0�b��Z���j���=�|���{��o����/)](;BￓP����bH7������qUWlz��!�!��{{}CÁm�{��v��۷����_��"�W�H���l��ϻp,�l�B�OA�p*t�F��k��g�#q���)`���GM�eh�M���>����b ��y^���m^̇~���� l���1�}
t�!�5!��������=�q�~��t	`{o"��u�0����O��E��=�p�sW�|D��}	��}���i��w�
8҉F�10t�f�g�nz����m��Z
���V݅���D0����d̀@	^W�Q阰q!����Ie��E�}���
�r�^��EO�ma'��P�ֶލL��(�t,,��R����>C{[�r=}{Ĕ�<�h��2���A������`��8���t!�xd�5L���S�ݧ1:v��y�0�������|�����Eug��(��s��*u�՜�	��`������ޘ('����i$��0I<z�i����@��8n�OY���&n�+���u��&��ٮ:䥫��!r �&���9C��
 �}��xe�G���S��.�w8��J�p^\�R�o=G�_-xJHR�,	%�7��V�aX6}|��q��hU�j2l~^���^��5|���~0�,�}���|ŕ�x�r:B4�0��7FH��Z��g`�^����L�׆;
��(pYQ�����mJ��M4ݔt�X~ˍR���S1�힙�,�3&wu��[��!	x{9��C��Q]���*�;���~G��?�`�`k�G�0��e �u��s��0 �$lɣ��8�<#ﳙ�����9�e�4��R87_$��O��"��],'@�,�� ��~ѵ�iC#>JEeeL�[m�GNC��:�}�S[�m�� �..g�lN��\/)m8iἢ��r�(�g%\�����0.Y��좸��S�T![��F���% _�Wd#�cIQ탴)>XZ��F��~���� ���F)�V�lS�ڦX�q'��х)��Ы(����dIm �a4�G)���󸙢�(=o#����g+���P4���^�z�����TЋ�/���}�f.ff�\�v[��������i�[*[R)x�寋[�9ap��ȥ��^)�T2��4b��G��Qbf����pz�T�o�?6�_�#�#{��j���̻>R'ޫH�0.|i�TD\��O�����/����_�w���C%U�}�{�{�g�WF���B�p%8{�ڡp/ߥ��}�ϪTfN����ʉ�x�j�&PgU1/���B�b1nB�9kr��e����9)��LLb�
w"���C^���ޗsƜ{[���=Q��.ﶋ`^����T���z錡�0�}r/��2m�o~���@��
V���vZj'�{4�&���n�3�#�ָ鉪$�[]�n�]+��H����	,g[���EBMW�d@E\�x���LY��K��`���7Z	t�I���y�j�8��(^￧4��q�W�{�J��#�> �IBȽ���_�o0�����%� �}����/(�W>+7Kϝ�-���K����K�%�<�έ�2����ϱr�]��	�Ό��}�����ȼ%@@Y�R<::�h~A�}�m��A�)D,�C��b�o��Q2���������L��r0b5��d'YG=��,�r�}��[�u~������A�Sv ���o��"��qIK֔��ޢ
�:1.|<�[���ϡk�I��]����+����<ou���	4����C���H��L��x��V^�˪s�?�oy��%%0��4�"1�B ��eP.��6�"�U��T-Uҫ����G1�ˎL���;����k=�h*��/�>�/ @��B�B��&�i��u���=@�m���؄��8��A�����,e&%#��������s��}�ŭ����KC��<���[V�iO��յ�����}���~����W(E�k�~�0 �*�R�z�?��P�(q�����?;j�3�T�4�0�b���x��,Rl�m�V(|@O���,�x����0"I'=��&@�.}��t�'f(���jP��65�5�I�xo�\	#�=wP�U�D��R��ס_�~�}�?S�%�M����e�hߏ��]9Q%�������+�l�dq%U#��6�p��u~	I����i�20A����ީf%�$�o�f�p���r�V��+"��Lڛ
8�F��Qn���2{�H�l���b�y�4-�:�r�J�� X�3�^��0;���͉�������ۧ}x8����Q���m:��h��>(kg��R�׼P�}|
�p'��f�1/\4�&&mE?�_�k&�>s��h�Ʈ�J�z�	�0�a��7ﲒ,���{��������ӛ�$�C�[�j��ދ/!4��'D����v��<��g1�>�;�X���a?ER��L|�,�3�R�aU*YSØ�����"��bVg�lR������[E*���LUe�10���_ޤ����e8pi������p��0[�����߱I7��Т>�S3G/����'b/ڒ}������6�],��_d�B0��b�A�b��'9��}:�",��[@X������!>�J���/*"VZ��D�����~��ƭ̒���j$���s���Gr!R�LX�W�e��Ά�	}�c���h���U��|�R�N̠�gA	z���.ض���E�N�Л_EL��h�I��2�;¢O�(q���������1	�q�vt�|^��e�%X������O7N>^
����/~�ymg�.���m��uǅ�-�L��:��&����(�"�ƶ����
�OeeX������`5ν䗊 �X��~V��+rǆ�(}��`f����5��Z�
6�1 �d�Mb������hu�?��;	�+�}�"��RL$�EHm�6Lm���>����'�9 Ë�4����tӣ}P���sx�a&���\s_���8�L��z�}6����ս\X ��(���A�����>��r_��È)Ѫ˵TS���H�@��[#D��������)��g��H����9��;��_?z���恸w���It������+b��6u��H?��� ��uCt1�������V�+L�l��n��=��LQf�U@7cTTԮhߩ��ㆷ��ިy�vʉ��F9ߙ�-EU�u�Z��eX��UO �8У� �^��S�*�ף�s�f��6o��y�L{qM�(^}���mdܧ�����c���@ 3V��rF`b


�Ќ�Ru��FʁB�4ܻ[��*�sDFBdO�xp�������/�n�S |��S��@�T�L�"���D���u��Z�ߪ�U�3e��~���E����H� ��}�4�'4-J�����hak+e��!͟8� S�ު귤��Y�a��'�����ޯɹV>����VlӍ�f�Obb���͞w��Ҝ��C�s���t��'�!�O����V����"��bٳ�`0�ȔI޽{�����Gr�N�7m���0%I�Fj쉽�Y�;��e�U`MG���p�H��������si�?��9*,al����"� �f*�������a�&��O$�u�` i��hd9>H�����Y-4�����\��6M��C�����'�-ˮ�cW�9B�O�n�D����Bf>�%{l.�3/;I��,;��/ckf��פ ��a��3U�W�4G&&b���dhW�=���7�2�ҥ��ec��Si��������>�`�t��f�;����!)�#`���HE���"�07��N7�A=E�Q�+���a�D୰��8[�Y �s���ڀ�Ѩ�z�N��u먀�UO/�O��RKars��!���5x�Zpc�����$Xg)wߪ�;���R4X�� ��W9O�o��+�!kF���b��Z�o��"Y�ݼ��>�ǜ'c�o�u�:�����gg�bk�����P��0��uS������o��k�t��f -�Y}����_[�;�ٞ�dI�q8N,*@w*aS"c���t��W������8q�	�d1�Ҍ1��8�`ݡ[���ڛ0�i6���BJ
�8~���?� A�ʲ�%���m!���%&���
�nF!w��X�����N3���?}�N���=���8.�/�SU�U����w/�Eoz���V�e�=:W��Ǝ���e��~�g�%��(��(݁:O��80����P��LfpU��Mp�S�[��ci)��W�n��Ϟ_�\����ך���DE�</�!hau�,,s���R��D�e	zC�Q:��t!��d��&�~�d��{(���Z�
��0H��KcɄj��(�c�Ĭ}Ji^�(��dP�G��w?�80����b�o��}��%�@CUM��\G7���'�.��b�,���Bw���=�e�XRCT�.���o�����z%�4�i�-@(��K�~���;��E����̻wy&��$���+�\e�K��3�V��>WD�l�U�2xx�!�K�-L����PUv�u�Z.��9��с��/��X����.On�K����g�$���D�����zz˼] 	r��6��s�i��H+�:(�j��C2wdtt�<Ņ��G�;;,�G�rA��2Ɛ���s%�&FmsQ��ym�����a��
c��͏HH&�����k��9ݝ�~��z���.�ƽ�N����oNP߼VP����v��4P#`��Q�w؀V~��ZYU�	>X<���D|W����Tqyq��$�iS��k�)'��	�{�-R�H�]+!��8Tkݿ~�g��\�f���<h{�5�Xqxv��[u�w����� j,�GQ��K�'�("&�<5�.��Ҭ�.\��	����%��,z�" 1?��,�������)�3_�'z1�Φm��_3Z$r�\��z��Ub��g�4E�� ��^�NII)��$)���]\Hb�D>����P*�}�Ւ�()��W�,t����������O�(��F�� �j1�º�FFElX���A�(�F�#��\+����`���b�q�VPG���E�s�#���=@��M�����g��ǲ��nR���v�q�~��=<!z��r���q��9 "g`�_iuj��~bu�˳�O���a[��V��\wm�$���
� >~q��hO|N�cc�p�'��-&���h�YF����1Q*�3�q��M�77 :���h��;��6Uذ�Vr:�&��PT�@�4lf~ۿ���:��){l��o j������xK�ۏ�v�C��ی�&���п��F����D��)P��h7B�72⪔iD�B��8�����[ �4�ЀH���n��O���座?�;t\x���K�\��q,YZ���b.��E�q	���� ���/���f�یwo�'�f�k,�j=�[L<^��9��L�b��t(}��}G��*wϭ�gF�]���O$1�T`_=Hh����b� �㮏�'N���Ϙ\��c�t(�R_�����r���43N_K9�gŌ��72���&&�(��s�?y �5!�q��rr��^���q� d��E�D�K�j�x�꽵�d�A�O΂�6��nz0��1aE|�3��H��1�������Bکok����י�-j�Y�M��qh�y��wi�A�l��3Ѻ�@V�,�Ͱ%r�J�kW�8e͇[S��;��O^�|8�����"�CK�pv�td|<z���V�{ґPP���u�<Ғ]�+qx�k�D�0����\(Z�Ĝ.9 �}�׹�d�WqՆ�@yj�d����C?��Q�x�>ؾ19 ������}���Q$gPI2��^�1�!���s}��f��,$/��"�I훣G�;�U,��dvr.za�Q�|3U�1y�Ty����R:���p����O*��vzꓥۋQ/jO@�*a�p8�_O�"C�'4`�N7��9�{䋪���V4�X��O��,R��`f�)��¡ӳ�Dh(�(�g^?�W�r�@��{?��r��)Q���D!��W�>'��=+��r�I��.�.C��r���>�G�^�Q&u�j���V�'OFFF�Ws�ŏP`�OOOqb�f�ɭ�}����_m�c��E����z�еo��﷮��~�K)>�6�iS�[����\�=�� �ê�vb�D���Z�+�vP�c���כ�d�q ���ٲE)�����^0�=�>���h�Hk�T';���&�y�� ��h�\ -�A
v�j�]����T� �W�����B�cp^���	���x��@�CyY�������4v@��w&0����{zc�~|g�GVo,3��XBݨf�C���n�;��A\|���F�0�<z@M����)b��~�Fz��q�f0��0b}���k#5y��X�E���'�\Y���sT��h)���B�X��j�N�᷊�����x��}
�wО���^ͻ�"�??�TRNz�����l�ׇ�#�q�F������U��a���`#	p���A�����)���|Y 5����, v44�X�Mw��8ҍ�}�}���Ĭ�������6��������:^��������_�$��֖�yԵA2�&�Lo9�L�Y%B��r[���F�|y3�8jo"����~�WV��^P�,,V���T����N�(-FĐ]�t�A��E6�`s��[�.B�+�DSH"~'�	X�t�n����Z���Q|x�P�1`�V��u��Ť|�EX�lqq����|���#�<`���*RC�.�X<�P�#���K�4ىFw"���[�����WNU2��K���w�x��?;�?�^�j�4F����s[9��b��mL��H���s�������X���c.��[��"1�{ν���g3o�:�:6&E�Cb7������2Co�m^8�����Yl�{~�����KgAش����*�����v5 ��d�!aX3s8R��=ȕ�D������r��m�ڨ��M��r7�S� ��Yaz�;i�W�kԵ�!lk����&4w�6Wu�[�+[��F�Ƣ�Rs�x 9l�1����}�M�l�6�G����m�?0���󁈍���nʡu��,@F�K��<���Z�� c�jk�_Ce��4!#����r^��;o!d���.G�'ΒJ#��E���ӧO���  N{��?����)�r�[�}^0q��AE���┽��-s�Qu�L�o��AoG��I���{�PӢ��K{��7�J�P�W����G�T�q6a�un�Z�@�Y]��X��&�M�-K�5�x��1��l_a��#��g����u�(��/���<��8�����3�5� *�����Q��`xu�8f�m�����z;�5����ܙO��m�%�-�v�������LX#B^DD��r�>�̍W_6Z#4H�z��/��H�'�\����W�{-��؜ͩ��80���i���=9�N3p�����Z�$IY<���WPX�7j���$��\zL$��-�����Aj
0�c�X%��B��>�Ψj�np���E���@�q!���ѳ�q��K�GzF�]���}@�t�TO�|����wb�^jx%�{'��WbV&���i����o��hk�'�OBo.)/��KT|���nnBB_�c86��9�d^�Ֆm5�D�5D����x�C��F������j���a �X��F܋ƥ�q�VVF��2���w����,n߷~V��؁��k���\���9��q��Z���@��z��ZQ��77C}x0K��z�T�F�ϗ�PW<f׻X��%5��7��~'�M�g��\g�K�@4A��-,����5�B�x�m�?[�(�[uhb������c@��J�t�`�(�����E�h8�c�X����-o�_���[$'g�s���	zt
�VVz<US2Z��KP�G�y�&�l^t����K�"�]uȻO����a@��/������(L���Rc:!��*\8�7�! i�z,��h9X���[4�l�3`�t�j��j�t$��:�8Y˂�D3��|�ѹ����"=�I�u��N��Ϳi~�G�������[�Tvq���SΚbsur���޵L�E����ScM����SԂq�A�	�>@*��b~�v�AUm��j�OP�w��[ R{𯨪�.h"��*�H*D>�s8n�������O� �|`W��\��ڎ#v�ة��;̖����]�oOB�k��3���>Ʈ��W�o��V�`����R]K^�6�ۊ��~��',�K�ǸI�2��
>x_/��E�ѥ�E������0�<4-��U�e����?��\��*�H8d��)�l&�8x��8�����"�q�7r�r�Xv�.��[�i׳ �v��w¶Ԗ�P� �1�t�2JF�M�@?���2v�:+�|��^w}���L���W7�DSr���J��5aGI��Vҏ����u<�L?a��é�iy�r�-��o*�)�ڳ��_~~��Dcc�3�������H��q���u>�c(m�Z��'�0� 2.�S<�s��^f���}ܩ^�=�o� -��CQ�ހ����(�NH�f������	W�;�bU�A�]ߪ.m5�SP`uu��i+�N\�1��;0Cn����Hp�� Ή}�Ƴ9�j_�����i�Y��c����^Q�jZ�uVs�����W�u1���J�����7�Q<��B��/׾�׫s���Q(D�W���:7���ҍ)�&x���0a�&�,�)��姱x�<�B���Zpz�9�1�������6���d~'{~�U7�=��Y?$��	�'VhC��;)>�f�bv���ˀ��� krf&R�=����dW�Z$��up��%6c����>�~p'yrO/z�-a0`�����q��ǌ���'_��skf�W���/������al�&2Re������Je��@�ʺ��!@�QJ!��M?�^l<#{o���{����4l�M8�vc��r�-�b��⊤e����
'DF�w�W'��	�h-����Q���ٱ�MXS�3[�I1�Q����T��MLL�Ӯc��eX����xpz�:���֡�?Ś�s�������^B�z�3/�KbYQ�K�%S\d�=���ǌ5�k^��]��+�{-��jR��l�:�'��(�btB���� 膱P�J�K���D�q�[�����|��;��x`�))߇	;B�J~�3�:ӭ�I��N��^/�bDQ ���H>ğ�E{$W����?չTҞ`�[���=���� ���]]r.� W޴/����98� ��/A��^x����q$EP�X��6γ�\��z�k]j��'�A���ҝ$/y��,�1őՅ�_�Y��K�=6��zha�rob�;H=�j�d�e�$����ez:�Z��;���Z��jO#�O̘��q���L�Wo�I�����y �/Nl.I
�"W�� @B�@�Ízj��d<���zc-�ϠfYU$.���jm�g����ʦ�4˭���9�	^�
�^���=���'�|�I���}l<7b�U��&�o���g��M=��<�u��s�G�Jn|z���Ez����<ر�Է�y_
�C�q�rso�Q�n����k�0��F#��'��
5�*���g����?~��-(Աw`S���1 ���[^J�3W%�c1!����|�K"��]+��W�34��{$�N�@��)���s|2'�O� �`:~2qw�Ta�ww��*��yV�����c��"��Y���Q���t��g��7
������Q�T�+۫5�o���e�n/�#+�*]��q6��8�|�4<��ETd��`�o���!��Ԯ{��J��))�&��H�G�'�����!bل>|P�Јx���q,�D��1ۢ�����u��~�V����	JL��Y �)� vi��j�����?�+O�C��y��ݰg��B�̥W_�v��\����B�[1��5��#�À4��Q�������x��������U5s���bp��e����ꘞ1�� x��α$��w�`v��A�8�,�&�7�7n���mW��Yd?Z�i�'�T&���-��������B+�������)؟�7D����p�*J?��������+��&/�Z��/����cM�C�$$�H�'=��+g��H=�S��^7���&p�P
?�>^�[����Wz�:g.��jk���`B{�$k��s�`�ƽ�f}_���^±�OfO�m�����,�	�`VHh0�E�%�e�AR`��V._F8�-#q��|�7��v(G\��T�cd��DM�ɘ`���J��ggP�22�s��y8�@�L��>���!���3뫧00��ǅh�$�GV||�)�>��m��U�^v���N�(�~�&���N?��׸�	#Q���R������Id���>z��^h�A��{@ez9�ч�2�h0����赠�b��Y�����4�x /�e��	���֝{��%�7!H��X�Jx����~'������"��L�M�ZF�m�������M��|6NM���N��^ƍ�/�c�kQ'�r�WWMnE$��c�|\-�d������m�����s�G7��W'h׌!g���u��Jd�ƞ�.�����W�oK�	���^��"���6/�(f�?����g�(O�+����pKi�&�x�^�&H���CI
1#,��]���.��H�;�ȕ�If�'� ����~�m�J��v�h����ѡ��(�G�t3�{�Og�I�
�Z��A���Nz�`��%ߊ���r�_�r���p=����w�;ʇ*��۷k^tI���~�[�����߬�#��?�T��v���%w�1�WWĬD{�F�c$1�����je�d�[�M�U25���&#�~�|g�Ķ�Ċ�B��U��g1��Z 0�*�c�'���>�x9�)}�&&}8�i�;}
Vy����T+ol�&�./�Z��33^[a�u�
����v��H�e�Q!ϊ7%�6��(2�׋�?�zpI�Xh��{���k�(I�G���,�>��_ĽO2<#�w�6�8�'���AW�7�dy�W�9{3���j�?�|��C�����j��R;��)� ����$:V��\�_C�-�T��Q=��͑��V��v��uE?���7�=�5F+�+ȗ2�'���iSTm���zN�,��$�A���Z�I0r����V7q��˽��D��{k�)��&Z(f���\`!-#V���\�;ρФNĖ�J�V�/24b��bD�k/�3��F���~��@-����%��~U��jwO~��9�n�۲/X�#F�AŻɂ�O�(����ֱp�~7�Ć���V�!C���;z)�t��R������*�OLMO?���n� (�"�<ƺ�}75*��Dw�M�1M�З!��x���Q�:۱�J��[����:#��(83Q�����Qg�4k��+�:��iL���h���x

$4#�5���.��j\�{H !��C���dS�)��$�v�G��݇z������a�v�v�O�vx	�O�qQZPc� @�P��<X_F>F$�vm<�>��6E3��.I9+��n�:��b��|~��4��{���dl��_��+H��Y�ݽ$��j5������_.��C�r�Cş3m�g?�/��3�@��9�X}��<}�׍��=$4HnE"���}z�}�e@�fEw�T��ɡ��P��/�R�XC}Z7���#EO���#q��K�Ě2�+�`\��֜��>��Ч�� �'M>f����D9��e��j��<�s���k��d9��0`��d��mEkC�P������b�3fXY��Ć!o=~H���(�'Ԓu��]�55�9�ZJ���p�
�f<����`}h�W
�y��s��D���#�V��<�
��rd3bp�8���� !i�D��5�^�	J��=�@�9TǳAu�R�G�b���~����7����g'�'zn��c�1�"�L�A��@�x�WcOlUc����}47���5E!�[w��K
����ء�M�Um�z=�C���cP��Q�Id�8��S ��C{��I��5�R *f�}aM�wK���������i���Yt��*"J��)ԩ8-Z��{QfXc��U��g��,�s{�<2�	դ��g��������>���/(v�e���<x�?���01�9��V�5-߳}m�R���+oR=�Bq��ԨsVO��W59ɀ�i�G�U/�$* ����h�}KѵC��շ��쩸�~&&=+줊U+Q(7.��(��s%�<�p�X��`�f�t���~�� �
?v�hKj�_<ZdoM�\� 0D�NP_t*���o~������h�}�N����u�2��	���[{B��s⭷�)�]��Ϸ;��c��$Z�V��Ld �A��BoTt�=��o�E7o��Ђ�ܫwv���kn���,���Z9�Q�^!ׯ_��c�h��+��@ƨ�B��i���������d��T��� �r](<(J�A�c�,�^���Z��.���� �Φ,U��T� ���5\�����g/���Z:����}��?C@5�~]��Y�����n�t���KV<��eAO>;����G�c���Mh��Y�P}�*�W^M�O���^�V��VN>���~"Q�m����6��~Ÿ�t�ܚ<1��#���d��'�p,��@|�#������!fQ'7�9�i-�C�\%�Ê|����������@���Q!�9�S�|"S��h�W��A8���P-&,'��0ǎ�:�eB���OT��(�����	�z*9�=B|Ntc�
��j��Rg8)�lZF��e��ܗU2�(��n�v<���Q>Q̖��>�.̥���I>*��lE�3JΕ�n�^F��>e�
eN3?<]�u�';0�li9E\]���Jl��,o?S�J�}k@���h�M��׊���<f~nn�w�|��~����D����j�E�02��k&u{G�GE)_������HGF6.�Ы����%Ŝa��daJ��Cr{j�/��fM�d&�����q}1˦���Ɵ��KZ�P����zB�I=���n�n��Ew�{-���زYX��'bK2�"�:�rh���[���ѿX�.}!_>  �$s��J��~^��m��-�^��Ǘ
��]�VY�DN�CL'�B�(���F��m���f�Q�,C1�w&ʠ����n>�������,!��|!TTZ�o�i�J:�w�B��6�&�u�Һ{u��ӽć9;ur�-=N����[�l���^��-Sd���߻C�� $Rt����M���Ԓ�g�?b�:p9�Z����x�%��?M+}+/�m�l���@ByT�1���ܨ�1�]2�((˼xV@קB��Z��.M����Ć��'Y�4=�;���-0�DN�����)`����s�Y}J�[�"�J�����ߦ��ٷBi�Ge���4J4>qRM J�������S�
����v����t)Ӗ0�W�g����xf~�\8�]&���c5���q�������E��9P´�(W��_e�i��ݧ��P�v���׋�c��P�2oQ�y��[F'7�џ���}�{w<�B[�oV(t��w_� }�c�x?�dI@f�E���-����d��ڏ�����n�#��($ʱ�m�b�/͎Q3_�%�� w1�x�NJ�A�'gg�����I66D����ř���b��gk��l���z=��o�����ӕ ���%m$c��z��~v���Y�Y�h<q[�F�-b��P��ƋQS���,��,X1��۹.�;��Y�Hmb���� ����6*`w`�)�q;D>�*�dWY�[�h�JP�'�)=�e���J�]���:��Fۺ�m!�����9r�4�υOE���|ۻ�[�~�����/`�Y(<������.&��ӻ�4�(��)�tL�B�v���3G�x*�ʮ@ā��#*����e�h���Xѵ���W��p�ʔc��y���N��?R�_�h:���W�^�����&��tЃ;�|��d��[�>�Wv�K�B�=!�б�+��ޖB�Dtc��d�~1vڔ4����q�\ɄZ!�P��P��C�C���vE܌����[�>��?�R�=u+�F���b��E<�i޷cyq���K�G��`EZ��Y�#�{'Bs=���)ؔ�H�ϚG�v����~U����ֿc)��8���#Aľ �ZD挵в,�>�-ጳ(��S\b���������c�;�8�s��O�>[7���	f��]�(-�;�4⥠��TV��
躃���V�кT���*�<�%!�rJ��kb��EZ4����8���L�y���>�?Q�;.���_��K������;k�~�t��q�����C�&t<�2��<^V{�w0��{s{n�u/�a1߫1/ #��?!H<��x�aL��%p��n����#n�~��64pB�Ğ��T%�� ?��H����Zq)��aPW&��ɭ���6͐�� ��]Ő*O��w����ߩs��J~q'pw!G����X�l���T���l�2v������CH�9��|�م<�h���'��c��*۫��~PnЩ8�\���u�Uvȯ��}l��溠;��j��Y��JLG���ø����T»�o��#lq��O����9�Q��v�<V�7�L���9��P��੠z�Uu���sʈ?v}�|H*��Q��lm$P��nO}�I��sEr�=tm<�(�97��~���>^�~b.[L�h~fkk��w�
�@4�62%��t;Zϡ��z3�S�Y~���&�*���-���ݐ�B/[�"`�?���3?��ayD��~��x��۵��j�X�Uĭ@>d�/�N��:Z�ˣ�̫�V�yR�K����!�+Mվ�)>>��G7*C���T@�$���񐸫��wI� R��n�͌�����rf�ga>ɠ�
�B�Y�f�7K��
G�n��\<A��Flx�Ť�nA�F�bڙ8��]�������!�'�q����}��U`S�Wx��آ�9X&-���<f1��րQO	>\'�����rbs
9�G�y�r/D�z���G�*���xĉ#ӌz4B)bv��l��}'�=<z���#��-�r[/>�m`�4��G�eQ��V�^��������)����S`��2,b����w,, �8h�;��r1靥ooݚ�J'�3A�My�fl���C�)T�Yq�ù�P�ڠ�8x���x}�]c훪�l�1��T�['��ߕ�z1��z&�<33D+��׷��2Z��`Te!�y��?�*:�����5d�4�6���I�Ige�ᐬ�܁,��(��c�,�����O�Hw�R�]��tw7Hww#R� �����"9�������#�������w����y�9�N��r18�e:�&�pZ���g�6�+B�ǟ�܄��:�+���^�޾�@K��+t��1U3lv`��D1��|����v"I��������W:}���QQL`�V�����H	\�WL��Q�%!Bs14�����n�_1:PD ����Ë'9��N�!��-<������/U�Ô�S�YBt�U÷9�JV�ɰ�$e��e���e���$��l�HGs5"��а�{��,�C�70��BaأL38t9(नm�e����__���o��&�� �~5�$g���'S�!Ǥh��1�����2S���� �i��ϔn���zO'��E���a�:�F�?^�B���Qn������XJ�T%�`�¢��C�!)B�L��J���RDEXkվ���3�0���lْ�w�3a��x�����y>���9*��E[�n0��0Is�!��̔���t*�����2B��0<*�P5BL�S�r5l�{��]kcu-Z]ƾX����O9���Y%��,�t�!��C���vߵ�h5+�*=�C��V@�I46�  �0c�$n�񶃥&	�,�$nT+�0ڶ0���s:+�� ��A��y#��?�@zrP�f�m_�۱����6��5vk�{n�?�Nu��|;���" ��(��X�a\��/xRZc8��d#�A��Kl�;p�(#%�Z2��|����鰐7�x����*v?���@�� �2�Z���q��Q�/�`�Jo�حX�U:����-D�ʙ�P^;7"�7p�ˍ��h�g0�%��%$��S=��j�͒��Vv�k��o�����y2�wiku�H�zF�A���_1���D�~󇳇��G��xbT\�����'�	��3��!���Q픝F�<]�ri���d��5�;n�]�<�t	>(�/��?v+���}~���|u�2Ξr�?�ޘ#�-��	��gI������K��xQ(�P��
�8(�1�di�xCt�s�n�>��iX�
<%/8d+fd+��(��2��q2�:�U��܈������R�:C����hT������LA�'F1Q� %�w��S�Efc90�gfS����}ϟ0�I��\l��0����`qN��M��f�i�O�zh#֭J�6�8�G^[H�1�1DB��ɵ��ř{~`a�y�Lу-Z,���F�b����i����H#`6?�7?`�r�qH���T�<�\1���匾�Y$"u'���&�ǵ [4�0�����W�)�H�($�����	��_�[5��Q1~nz����@^���O�B�>87o������~��*�jug����H\�9�x®��Co|r�:����?A0�9�P��!��J0Vo�EBԩDб��D���L��!sܻz��Ǽ���v��!ߺ|s��R:N�;d�(`�,`�C�)g���+ju�L��!�L�5�22�0G��c�v���ʧ*M�mU����d���a:����� ^l���r��w¹]?!R�G"����~/Lvqh����*-�~R�EI��R�Z�)x��5�]����,�X�
Q���\.����L�G�H����{~O��N��öiRUJ�M�r�o���۲����A��0]�w�7����짎h$�]VV!/Q��篿&�U�Hz48��֍{���	WH����	)u|�^��L���3H��lk�d%��;�ʛ��]�����zG�l���S�}�itӹ2WUd�]���I��d5*��)�O��	�"�d6�0�#��m1;߶��%!��q���[@�4��%cf�Q�G�I����i:6�-in���V9���3�SC zZ���e�Iϙ j� +L��zH�5��G��X���EmӔա�s�-.�����:S����������� �iBJQ�x�
�����|NɈ��]�Y_�`yϣ�X���E\�j������,�#�}��vп�gI",�=I�c���`u�O�L��x=�q,��ʔ�����8(@�yb��g<[��ԣ���{-��~�p�͔uR�\��\�a�*�\�0��B��__!d�#o>���0��r��q�����D���k����&ѫ�S/
x�[��<��2;,�]�b�L'[P��4B�g�C{�?���6�G�3'5.݋x��"�)��b�{w��ٵi�@U��9�KJ�7V���+BM���I�Z$O��Ó�Lg�v��X|���"0� F�'O�n'��AX�����/�)�����`�E���b�e��;�	�N�S��q-F҉s1�}F%��'/�+u�A����[C�MЭ�BZ��Kz#N�qm@ǆ��F�����?�?��lwJ�`)�9�|c��>H}\�C�ȸ���r!��|?�Fp.�+�~���ǡ�sr��9:�В/&����CQ��|ۖ��A���ӡ�֛������!�o�(��`\>�K�hx�v��������m��c#�����T��'d������Qe�@<��Q,-?�NT��t��|��<eQ۱�����O(�ù��Խ��A,��A�d�ݒ0���>��\X��I�>q9����a��s-�]��>�ߜ��	 =���ه����7{TD �~ԯ�F�>�,
t��)��ί�2B�W�cóf��Ko�Mr�8�y�;��N7&`N��)eH.��c!8��~M�	�6S���2	��wU?���k��Rj�W
���k�����@U+F��hn^���� ������W?���VJ .�ґ�!>-G��g� ��7���->���9'3�#Z�����s������a1H�hl�z�^��L�^��d}��I�/�������^�l��ò��_�r�WP�g�M�εujn[�Z��J�����{m��\����d�7��*4!�o�iG%�3b�Շ?�F�qZ�c���*�$�rՐr�~0pq�ؐ�,�m�{��>q����5a/r�K��
Ӓ7��鐷���-<��uޛ:m�γ���J��;Wt{E2��|rU@:�,_��)"�YJ�>S���>E���&R����+�ۻa�(��S�+�\�}��߸���y�6����o��%`r�i��5�^�94���� �����k��^x㿶������S	���JB�~h~oTa����ߘ�rԀ|�����? �����7��Ch��Ͽ��ߜ����d�{��X��1��wē�����P������h�+��ZL�\$�Ն
V"쓰D7��X�����p�n���k�8t���F�:*�: ���b��j�Ԃ����5�b�\��_�y���׃�:H��]�}�F.dm(��߲=E�8U�{��pԐ���Ó�5eZ,o����k	 v6|3�(�$Kn?�PS'���s� Kx�
�m�`@&�%Wwq ��',Y7P�5�>t�`a�����$�ԅs�M�3"T�����˼�yToА�\6�$�e<q~�Re�6U�1ִ�M��s>@^n�Dr��Y�G䐓�  ֙����%�YJ�;�2��w��d$�=�Wu�-�U9�a�/*7�&��N�_�;�u�"-h����DCt��bc{7Sʫ{�4a��!~�3�����N��9�슎��o��E��g��Ц#�2^2f>�I���e�յ#A��c������䎿B^��D�Y�c#*S�*?���|��RVml �-�:��=���a�M�*M������F5������������5��������ߋj��r4�)����\Ⴟ&=�\�8R�l�b1���C�ox�ҽ�&���)aG�U�>��W�J�=�v@W���(+�.���CઆW1�i"����E݌C�Z;B&���/n
�� �-Q�NX.i����%¡����헰��� ��� Գ����n�P���zߣfn,P&�.feE���|z>�~��f�M��2��>�U��cĩb�������|!�>z��-�%wH�w��p7��F�ᝊ��Q��JFA�כ����N��y7cX
�K�0��pR���w��\oW��O��R�	r���i�ԏ�؛��k>���9�c���d�a�^E�s����B)n�8I�t-��:
ȟ���&u���r�-��*���
��;�)�Ƈii~��,�� �GqD7U���Xû�N�l��:�oc��	i%���K��s�W�(UKk�L ��MlDCp����*��cG7�����CN�G#.TA>���2�����/Ty[��;����K!�PU���y��P?��¾�ƥ�~����ss����E��9r����N�yd�0�}���t~n���c�?�*ȍ������_�.'�"<�=����\���F!/yZ�*���U{�*t,��vYsv�Fn9o�M��������Ãk��qQ6�I������7��M73=UM���{���Hu��A (�T�b�� � ������R�&�)��0_n��x7���za��d$��q�Ԟ(����;�����ǃoW��&�	A�ikvFT��8��K�����HE��a�cݥb�3���_3�a����.S}g_���"[<J��^X�d����M��	 ���N�������bu�1�?ɂ+Ⲿ �e
��.���*T�e����z�:�p2[�Prg>	��01�Mt�aa�8�UhwaqG�;wҠ�-}�R�r��� C��	D�{{ �u����G����D⫪M��aA��������A�<q4���Fx����y�s~s��ّIu$���{O�6�V���-4�X�tPu��gqM�{�Ԫ�m�!٩������4��-w���p}�E�;e�����L?\�[!�����۞�U��[>G�q�E�$��؈�?���;�0�����Hl0~Yگ�8\b�ٌǳ�v6D��sJ�7���D�q��=����qW@��.R�A��6�2<y�M��_��[W����x����M�9}�B��[)��9w����5 ��`n;���|b�박
!�To�S���`2���Ut!����3�� ��x)��k^�����N���b]>E��� �Я3{	08e����d5��B����Q�iZ��l���!��`�2$�x�*��+_��t�M�e�t>�QZT*�j:���r�Ʈ�~j�G�ģ+����1����$x���a��Ỷ�t�'^$a���r�A4��������):�Y��ý��D�͑��n ��g�U9Ķ4�C7���&���H��Y@�Lv��8��y��2������:���͍�N|[l��o�P��KQ�*��A�\ Y�9���Xy�D��{������܎0�O5��A�F߃�I�73��~�m̶W��03��g�N�7O��.2F9W��m<�X~|�)PG���4�18JFA�U�n�.C�~zc��q'��L����R���O����L?�����R���"���Z�����A� �������f�ޔ�r���� xGXAygs��|��~�|Y�Jp�0����c2����}�A�B1��y��<B/���������֞���dIo�J�� r��:�i]����>)gX~h��#��Љ@=@�;G.i}C"�,��3��[��?ϻ��Pܗ�]A����~�/5��WoG��<����`9+P��s1�	�܄I���д�ۢ��m��N���F�pt�?��I�#U.j ��'
q^@�?��ߜ�l�uS�ߪ�;�խ����$޾��h �{7b�]������lݷ��#�ly10H�k������2��O/�G�,H���To����k>QQJ9 ���ɽ;Oq�4�oBL��Fku��L�vgW�~�#�R`��K�ayoJ���&��j�Ow�K���h��6����m%�_y�5 ���{ǫ\ԃ�;��������ͫ��>��� :���J-��t��v4�`��Z�76�������jM� 0ʓO^�����g�[>{<�$�F�I�`?�(�_���Q�����Ȃ�#R��?����Su+/�BZ	v��M���=�/�r�ڂ��0�-�a��)��- ��߂���xpAN�]�����P8Ғnag�Eҝ��AAKA"�E������;��n�/���.�ŵ��D瓀6�|�L�I�"����(&����}�Yf?9m�v���O�)���8�ٜʰk,/�8 �t�xMH����N;)@4��dܵ��%�X7�6A����HFFi ,��V�k��`_F�oʁPE��셐d�OlLw���S?��1�3�~��O*�}n{|�� ��;-�P�d?{´~�W��S���O��&]?��0�:����a�}Gߴ�2���.x��ŷI{�x-�'〷g�/�51tB�&2}���N��+s�m���!R�u�4���R�X������I R-^��������L?����L �˯���I!�d��E!=6���@����rk�¸�2��u�QXT(/�׿�_ڰ�(��7�+�e��������G#��+Ĕ��[��\7oo�-�M�S�p���C	J�-�A�}҆GaT����D=��79�]?�,g�#���,�v�G+L�;f��u&��u��M밭���7� q�ٴ�Ү�ϭ���>�1.%����wd�6��`$�N��B�k�Z���K+A|�Kd]� /��Ϙ�X��O�9�����x��@5<�g��|���/{n�Mf���Ӱ�[�)�:x1�:Ǜ�%�c��p�'Y� 5������xwz5�jN!�Jk{�V\�a2�����%���MQM�24C���qMXR�wP+����`���Կ�c�SKl���R��ʜ"��R��q���ִnʀm�?����o�gc��͉'=��^5�$�h$�f�#��+"�������|���dj�y���<���r�g%���@q�_��>X��K�i�,e��i�웦��5(5QQ��ϯ������m�PΆ����Lt�,�	i�� �pg�����,
��YLvu��<��$�U2��1�K�:i8u�� ��cA�<x�T{xu�-��V�{g�
�7�L�J��x�ߎ������^���PW��]\�r��Z �w��fc�ނ���VE��;ʡ[p�&tb),�C��7C�v�f��C��U(���P�vqZk։A���yçc�C�Z�1���)�T��18�6�$�
Z^�z�f2h�'cP�8�!��~W j= ���c%��ni�6 ��D��ѳp4k-�1���Q���
'"�:^�J>I����LTċr�8��`b�bC6�o��8���5����#���;L����=�@��w�w�1���aҭ!Oj�|�=
������0�2�>�J� �,w=��t���Ipp�+����׫��bv5����#���Ի�b57�#�m�P8p�Q&��TGM�X �vɥ}O�f��?��d�z]N����9�ܷ"�HI+���%7�t��r&=�k��ߒ0�K�ӿ���'4�?ֹ��mL-,�ుi%Q���6a���3�u�)]�ݕ�U�L�")�u�y���IW����Q2b�/�"��Yfr�/vP��>�|����D�6��Tj�Q�lpL�o4��Q���ݜ�z��=[��e�c������Xu������� X���2׎�M2���V˓�R��ŉ�&�'� c�?3vVb��A^S�����EJ<i@e<�ő�β���cg�x2��7R!�W*~B���U?�����ZF�_Gx�4�y5�z�_������T>Y9��=���s�����(��u?'���A�/�F����!�S�H�����a��1��M���U��a�ٗVl!���ʋ|���φY�M���
ȇE�H��-NBĿ�+VC�P���g� �'�s�g.y����tM�~� "�Q�Ar<Hv'��E��p�n�*¡��w���⯮�R �?=��8и�&��gK���2��=R��|��K�KJ���_ŻVlS�_���!.����U�j05���q�� �����g�)��ۭ�˧r^=A����ro-��-*�m}�}���7̲�=A���P�S�W���e)�7�����^����ک�B}6�#��s��Wܷ����[�߼j�$Q�&iez|+���f�$,Y
X^7c ���D\��k��7e밀-��X�0�H��.�q
�������/k-'���{י����T��D������N/���X�Գ�����Tg�<8`⥄<r!GC��U��ؤE@��*O2\�{:x�������L���+KY �"!͒S�3V�K?s+ ��6<��ʀQ�Bݕ�2RZR3���{��AIpe�ş�r�L1�� ����-�~��Z�'+�M���|�社���/��kⶱĈ����\����Ƣ5p���uR���x+�� �Ҍr�r�'��v�n�t�l%Z���64��E�T1oDC�4������om]�Y���͒L��]��g�38NJk��J��̄"��]ȼT��|�\�s�������Ỵ/�4��$��
ʈ�X�aZ2v:�����Jfp�Qf�C�z����	���R�ƟU�KP�;WQ[�������� ���:ܭqh=�4U|��(�r�{����&�{���L�&��(uF���&C/D\y�6�U�� ���g�X+L���z���᭒��hVٵ��Ac0�p����x����1U�l.��֠�?K��@��39�0gn�W&s@6����6c����@�G'b�m,4{��`[��V��zO�R�]O���N+��K�<U!�)CP�h
iN�-�f�c�Km������j�}:�������HS&�z=UTX\��A�n��Vcdxqw�;�㨋i;��S����%���������	�*�K�M��P��ˀ��突��;��w�o%$���\@~�|\����DD��r�_ُ}f��6� `��i�*ve�P�H�U�2��t�*	�} ��^4[�f��X�q|�3��$�c`����f����o&dw�M���p�7��:��Է'��J{�W�ߧ�ܝٟ�A!�Sk�d�K�|����6�U]�_�w�W�#�f�a���Nrv_���@34�1�N�q��q�H���i�2n�T�;� ��_��'ǻ!�Z[5��.�짋_AG��uM]�'Ĺj;3˖M.n�������
��9iH�v7�8���S�k/�ݪ
3ȫ!\V�ɺ
�3���2W ��88�Y�
�q����y�$x�ĂFfg�=K���G������ޫQ{{��E�ᄎ��_,�͛NM*�[�P��
s^��V��'*Av�w>?�![���8���!�P1�v�$&�=|-��.�������J����k(5,m�:�A� d��@�f�j4iZ�ܽJ�p�73cc��|::�!؋߱Ws�E��ǋ�c���mһ����TΈ�2<$H�d��soW�0��	n H���!��7G����ƴ�8��>>��7������kXką^��U�!��Gw_X;O7��\Մ�j�J ����5��U�Ѳ?��oD�s!}^����^�_����$�L�^�����i%P��F� C�+��|\�ZJ$c&��n���9]H�V��A=DӸ�D
:����WBi)���+_"�u�&81c�#�l��CKumb����m58]
ǐAi_=��8�v �o4��T��f~��T��a�=NXVf���_��a���򚻖���QHb���fw�g���a��Q\��씝�Uj�2�l
b�>�Mv�u���f��o|�_����W��h
p��&�Y:.`�Ba�l�	����p�����l�` ~R@�x�i��,���Jg�Yr�ҕ�������#�p�	��؏�J�2����m0�,r�~"��oC�b�$�Oic�
{C2������Ex���6_ԉt:_�/��NA�jiο��D�2�������"�v�!�S16�C�ۯ�q�S���9�Rߍ �]��T��ء���r�os�9o��
��#@�Z�r\��>Z�K�@Oݬ��$��{9�V~Z�e�W~����N7����9��r��?#�s!:g��������L�Z!`gE4�x�)\� �V�Y�Ò�&���~�����.�1U�Yq����\@��en�ln/��%�/~���0M8�r�4FB7��xG+$F4i�=��yMM
�;f����z�@������ ��׭�4�H������Ͼ*��w�^���ى�@�!���W� �=�N�����J�m*����b/�������������n�t�PH�<d�wN�s�%!�F�=��P*�\�kU|���L�3�h�R�)���P`��:�#+>U����">Z";��\[Ge��ư;b8V�-/o��5��e���l��籫�9��� �yS:e\
I���PJ�G��­��C�3�V}a��b*a@�.�~�x�Q�k�m�1d�7%�P��ܕ��>�����,��� K鮛fnG���_(���B�_]W�>�S����ŏ����s��6]��OZ��5���z�Օ���,�����`<T��gl�Df�|j��$�W�.{3.�^	 �b��CT��E(-=�l\�(؅b_���	�^ޝJ�@����Kzh-�w�� d�����I3�����6`��lp,5߃�����g_&�6C�
1!��M�ض�^��`�`��O8���'ݮ�䊳f��-�.<F�^@u�[=W!�~���b�'^��:��b���{.�ϝ��o�w�o��>��eg�z�����Z�Ð�=�ݧK�o/�2��S����v��7��;��[U�V�#HT�a�O�~Ũ�-����$���R����Z>:Xv'r����n�)
�uA�^��/� �zl9xn���p��G17$=���~�y{z�f�G�Գ�ij0�kթ	K�}'�z�;\Z��.�쏰e�d!-Բ_憣���6֦������%���0��	��  ���f�螮�1��Gt h�&h�nx��ح�7}y�Ve-��ϼBTs(����Z�1)�
x���t�����{ғ�Áiux/bR88�F![8�#�*���������� |Ej�N���ܾ�Q�'EuP����(�a��z�b��.��@�|\w�a��9���{�吊�VS���������3B�����7�}�8��2#�P@/2�c	��u�ɭ+UVD X����˽��� p���>��܀<�^����`�]����)����ym�{�S�Bj%��&��en�åĿN��G�@���4���P<�}a�Ȏ�?�����<:����_�E�V�T��Pd|�y�����n�f��r�[D��@#�sH�ܗ]ǉn݊�,L|����ѪcLD�ڸP2*��!�jۡ�W'��z�S��w�Iq"O��I�<�(�C#bp��/h�dv"���MP����)���f۹%c��-��X�q�L��𺝫���$����?4��*��S���Ќ����g3�}?�_M�~�6(|�1L)�`�\٥w$Ү%u/�=	�x�(�@�������n~���
���qj�qWBZI��ѷ�zG����Z�6^P3/x%|E�r����f����������v�mЉ�,@�M/���Z�a���؆Ǻ�Xnn��-7yKul�]o��^�?���p����ܽ\�3��S�����gI�s�O:$��6\Ȓ��#��n*{�wfbL؋;e��]���v�s�\�Sk����.�?��R�Ĉ�5�͚�\�����ƙ�ar]� �yc}-:�C���o���J=�F���o���x�&��j���6�F�N�.��uR�#o1�,]��Y���r���4����`K˚�<��S��BM����zo�N�[E��.E6��X:�2�#�N��hg��!�G/@�����w�+��#�Y;x����ؚ��VU������!-�	�u&�Ƅ�`�j�F�N�ӷ�"�Y4���Kt�z3�q���q��?M?�����=U:�Uw_��ERA:��np�E�d����kK7Q�m��=���$�*��Z%|e+��߻o��`o*�1�g�(T.�V��m�����w��^7d���u�W��%����`���M|���k =�����;�����������Kz�����<R�E����N�|N�mjW��u�~UP��\'Χ�h^�1�5[��r�������;���bo���jxG}��u�֣f�6��Xn���a��'ܹ�3��/ex�����:���w{O�2ϛ��k����Ҵ��pL��� ��*��m�T��V�<Usb�3|�
/ճ�+��'P��<�A=A:�O�j�O�XP���?���di)�y�#�3TB%>�	~�u_�V��!�ʎ�M�h�@C8;S�LV�V�mA��Dr�KnQ�/�aZ��!]KD{v�&˖���t��`I&4.�W��@MLӸ^69,����G�n��2�~;O��4�yU=�TP��3���mD��/��h3YQ�53�Z�ɢ#6p�6���8kAC��	Q*�U�=����ю�*+#��nR�5ҡ?��K�QQ�`�N�����8���U�����@�^�Z\�k��\P_�O@\�e6O<>�{N���^���-[z�yVj�Gv�k�{����j��ǒ�]\�:�'�Bd�s��B��&��w:��o/��PSL��W���V�-�[�n��m8w��u���\�_�o�rb�]]����9���~�K<�E�B�)�A�X��Cp�zO~���a��Qf�!���.; �0	�!l�����r��d�t�1i�x��|j��Lm8|S�no���Xf;�yԭSV[.�n��N�B9�&cѶ�x>Ѷ!�%��!�\���C$�g�6>ھ����Ϛ_�����o/��$����7���wW���-y���G߁H>52�����:��p�k@���s�H����|Y���1][�q>��49?�F���<����E�>k�r	���U����n���8:H6l���fLa�g��X�T�"E�ѳ�}w������^�H_j�'����=5}O���5x���Iʹ]������1�.�U�q>�"�;�9�{��s���I��^.xָ)P;��z�k��?�ͣ��IGfX�f �ߞ�u�&�ת�=�X�"}��#+���Z"�Z�Α?��_'�����pȞc~ӛ��q0Y����Uw�q`����=h���������ϢtD`v��&�_�V�!��b�=�!T,���P��3�}a�>已���2�r�K��Z3��==�]ɫjĐ�h�Mx�8[�HR��H�ʸom
ycZn�\��K~��!D�H{������������l٨k*S��Y_�M������v�z�b�$B�6�Y{�cи�4}Ά>�G���z>�Y���1
f'�y1l&���S�(Z�W�
���T 3���ze0�Ns<�V�S�ʄ(�ZG�F/�q-�n�?��3��Z���F���E����D�J]+���M�w~?=�B}u�����.�ʫ�i���֞Vo]�1Ek�>]���8:��J]_9��Ox����N�j`j��"6�2@�@ET�c]n�2�6Յ��t����ה�]��Hs|�p~)��AK4�Eb�gC;�s��AZLϾ�k�d!��f.Qz������Vl&gDa:��3�Ԉ
���z!#8��Z���A`�BE��4"�g�T�`�M�H&�.X��-Q����p���+o�(0��w�{A�_���𝐗ZPo���
e�W�O;��^���DҶ>��m��I����E&��_;nJ2򦨚�;��C@*�zf��-���n�FX�XƘ�r��3��S����T��@��p8|�(sf���z��	D�Uv���إ5C�NV!E�<���N�KWp�u_����E�R��������L�D�]����m��?#�3��%(�IX�Ԩ炊$�5R>D�A}֢�Ϻf���1���@�!�WY��4E|��o�|!�=��)��t��S�z`�����W�&B���J{V-=^���o���j,Q>5�"7�2�:�M���G�i��13�{	��M�g�36!
W�&	�1?��M��EC�M�V]��o�-�:ߦN"y\�%���z5���;Q+}/qO�����a鈍r���ڗ�מ�Y[͝`m�����3f�.�h&��9
&4��0��|=��BNhZ��͑�r%6c��ׄk .��꯳�W(J���!5[��bꚜJ�e���^X#�jN��س���(�PI�$�� �*(|y�����(Zt���짷RɆ��a����]��y������KB���UX�������1�(m]���;+��8�ߚYK��M9"LP���CB��5d�jh��Z1Ҵ�+�U2�����[����ā�:#�8�.��۰Vʂx7��+�н os��Y9t��r5'��(�����Nӝ���	�����'�%^,^�&e\�?*��Z�ZAU'4\9������1
��E\����'���{x�d��(�Z�z�MA^�v�d����0�F\����M��9S��8��r��aߞ<��$iE��{a"��e2�k��3�QEW�$"��b���_'>�[eT{�Ӯ��J[�<%.#�q�㕊��e�����D����`��>��m�g��Ѽ�T�/ǒ6���Þu�1���=�\1�E[!F��
i��b��Â��p��1w�r��LZ��=�`Ro~�EOzg��DV~�[~89�ð�[?�w��?��|G=���rf�̆W٠D�뾏i�7�R�;�i�O�ܬ�v�E�T��g�mM�Ⱶ�ݷY���CF�`�
D�olw����;�q2x{���hhڟ�^})�:��v��ε�J��ܸV4�8?����qf'ё˅b"#�$�&�Ϋ��n}xK�i�����4b���D�#z��GKV�ۑ?�[.�J�������D`�W^
�;���(L�n�0Ϸ��QK_^�Kg�ː�Qހ�q�N��QP��(��b�'z���n|��>�
�S�y*���!�|@��?AE�\�99_�L9X�o�E��.���������� �W�"c�ꯦda(EF%K�qӣ%�("���v|��ެ1k[z��$���Hm6�p�*�e��&M�	�:�v:���٠����g�P�mg����&��� ���K R��N֧�����G�C�
��l1�H�_�gEUN�lf���Q��F��l��R�7��z�4^��?��<�iòmj�� T�1� z�_A{m�C�Y�D��ؕ��ѩ흞o���SUoKK���Q��=�O�U��k�_�_ 3W��-���<_�o��j�D��vN&��iL=����^ U+�����J�FKd"٪�b�K� �D'(c#���vpE�w
([�E�R}����cw��b�#�j9_��^��� ��)�| �8�����;�yКmn�o�y�9Iagݒ���|��a=g�|w(�"����7f�9��e��g�(5NCF5uz����E���+�Ն'0����^�th]���$
T�.rs��Y�}|rƳGu�iZ��:��wH&r`dT@�� �{�*�ޭ��4���K���[����0-�De��W�KO��h����/���pd�xB���@qmQ����"���	cɶ���p��̮�]���,p��"o��Cߔc�8�~��!d]U�e����]r���� �%OP-�(��EF+0uW*�u�Aw�Y��ހ�yV�U�K�bL��c#�Lhvv��g�P�A�n,Toc,��=}�O)q��k[�U��z��C���OR�/���"UqO^�Ր������t��"��	��/�ʝjʙ�?���-&�͋E�>�s�PZ#��VN�t@��+>:3�WA}�����R�j��{��э�Z�n7������lk�Y�~TrW�!�hɁ��Y2�ZI��-EB2+��н�a��0լ�*+[v������ϷW^hP
�:ޯ�M�Ry31�ꇫ���K��ߜ/���	��Giy��G�A9��U���Mx#p�ڑ�e��Ԯf�G`hg�E�MT�ty߾Q���v(̕i����������~stp;�(��)U�3��'J��1�?�N/�i|��$�>�	(	a),�38�tqᢲ��Q�0�-{N֬ڤ���ݶ�d��h�$%��z���U���jMl��G�"P;gL�l���'xW��~��,G�M�o��T������s٧���$ľ�i�	x����ʝo�¤���Z���o=��e}�<B�i�+�tG}5� =�q�q�K�K�~J�$�%נ�����`��h�4�+����޼�8�˦D�q��7��֤�l��h�~�S���Ay"��P~�n�=���������^ �-��b�f���b�3 �%T�x��S���Y���S B~����/�萔ֺ�U����[(:E����'�(�l��op�O�{�;܏�uǗ��#�`�!_=B�Cv}
�+^5Ƞ_a�*&�o��$��F�~�#@F�����O2�.��x�!hē�F[Gy�6�`#R����y�z�j��=���3I�����x�`��!�r��{���G1���&qB�'4^�6e��Z�#"��W ����Y|Vy�3�� �(�%� 2�*��%z�
�H#�&km��Ƒ��ƭ��[C=T����$�:~bX�Nՙ���^t����})F�cq֤�V����t��d��Hc�(��������4*���>f���g��{�y*_9  e[,hc�h����y�|U#~Ԇ����.�w?9�{�x$�U��Bi<�.����ۗ���O��o�G}���jri���u�}����kd0��P��$^5=��F��|�)4HL���:+d%�����|�D�^�0?�Q�8M�Ng�1D�|Y*a��k����]ƿ�W2�;�8��"s19��~̊�����8��b���^�t�*]��{ˮ:�-\	����%8$�[pw������!8www����������'�`��U5�#�f��S	�lw`�{��8�&�;�̍K�TR�)���:��!��A��<�~DWW)
��Fr��,�e����aE�Ph͒I�d�N/c���O�9C�\fh�'qw�W�!������Y$F��0�0�nD#��S�8����ˁq=ģ�p�ˎ��n6cG`�*\I��ûGsr��O�3x��Π�Y>H_&�I�Z��^]�u�EQۄ��U��,6+�4�Rf�,bأ:6B���ϮҖMfmn^��^BVsI)�(��E0����i�7�K�L��Pӆ��)���\��I�W��3��)핰藦�?{��Ί[ �q	G�A�.ӣ�E#��x@�����̹�ƙ����I���Vy��ϯ%X���V|�h�^��^�b�_c�bNLk��{r�}�x; 6O������^��JHk.Bgj��p���g��:r�g�&)�V
�¾��2�L��v�i�"�	�S#��v8Xnc���������+?��MQ�.�6�(B�R�|��MƆ(�5.s1ws�5�r��0-�fap����,�0�q�����DV�I�����'�KYsY�� L ����R��JC���f�v�|y���u�hE�3�\��27���� e�p�]�W�Qm�bN��8d�MNqf��\#��*H3����r)`����Xrp�΃��D�-����?փ:]h����/���4�jk8M��G��,�iц���A"8�pt����/�!~ز�\Q}���#��h��6|I�fX�T��ۍz�Ѧm�#��؃�<kb���]�LZ�6�,����}�-d�9xk��~ >/sșMP��x�7z"��RN�PF�Ϸ��v6�/nۘ/nM�>���=~��gm�>݈�
�����oue��y�_z���t�O��O�	j4��"�$�?>�Duv#�͈�5%�=�3e��Mͼ���?����wl�Ce�[i-�<�b�"gM�2�6��d�J����>�!ǎ���b�d�I`͂n�]Q��Hvc��k�~JGM*�[�����A������Db�$�j�.s���j1������ʅ�h��2#��&�	���m[���-?�c������k��b
�yl'�4m*.�j�[R�h���i�0��#���:w<�T�Z�Z����hZ��� q�O[�Sh�$b��*V|�?���:�g#H�{�<a��➠@K�����Z� 0�k8l<H|�+Wd��^<��#�0(�u���o�3N:Bšc'��pW���]�mE�bݡ�$V�4��]�k >�t�oB��el�˶��t�n���:9"\�,<1��a�Bk�����E���g.¶:���oӜ.mC�*.��4����a��Kq��J�.]W~��!\��\��ወ�t]?��r-�O�V&e�[��%H��}���CIK����L�Ro�F�����X�G]�'��!c�{hr�f̯,VR�|Y�p�.����|Jv�A����T����ѵ��c����2X�'4�?��D�YR#Agbq^��	ޢ;D�r�G�ó��o������ߝ�h�����~WF8�K�-�܏���ֵ���<�}�C��w�����P��#�]am��E�ݣ�3\|�v1V���� �w6��j�(/kx��aJ����J��W!�Tu�@?ΡQi�%�����	�/�k��^͈^S-a'��S��B��F���x���_O5�u�i	$鈋�6y%��e��2�7��Y��\�ʶR��n����u� ��1E��reE�a;e��8�� �A��_�Z���<:3f*�tT벡'�9�=.S� �ųUY�5��a�ݸ�O�0�K��V���7�`sdw�dÓ!H�'[v���;��9�,�!m�7Y1 ���9Ӝ"�6��M�329pbZl�ISQ���]���d�T����B\�_xTh���y�ah�Ħ:�K��
�{�����B��*�A�#�j]	5������Fꘕ��c�l@%	����|�ɋ{!�R�e+vq����ᔚ�P��-���rM5����"��wn�H��l�r��?	�AC�9}̘k[݅�M@�G;M�=C+2^�YB3\��p�W����C�o{����
/~�ן5�?��!�U�0��/Jm6հ��)��6;���Y�~Ű�ҭ�������I��`B�aH�V�`n������C_+<��"`|f�7`WKt�E��mtX��a�Hh�7��B�l�����J���7�#�RT͓�Pb�b����9C��R�C�fT��Y��lDu�����"�Su�uH_;��]0�y\s9�����ѝ']���gU��#��.�.�"f2-�u��iN�.��e��m���%�oP!G>i�CŘ�5P*����yY��S���sP� $1�lԫvK���W���E�W�-@a���ޭ7��Ђu��ex��h闤~������«٬G��'��Q�ʯ�]�2�ymv#T�=ϧ|�AZ�|��<�����?(ȥБ���o�Z�<��3�و� j���H�e
g�,K٪�w?��l�,C�r�~���hrV�I�/�}wBJ,�A�O��:�Wa��P)�Ϊjʬ/����s�n�1�W�Z���Pl�9�id�C��rײ�����簃k3�@�aK�Κ����q��9� Y�}�o�����~MA�$A�D�֧�E���<5�B����kֳ0��VK�9�	q���?�c��s �hǑ���M5��8�Q5�w��X�d�A��.̮ht
#�����T9?0O��ui�O�6b�?P���>xȊ��7@v�j�~�	癮�%��rհ�Ea�ǮE���tV�k��QkM�DQ�\#����I������N��0��ӏfbQB��K��:h>�ؖ��GD�.�ߋ}o:=����M̕�N����O����]B�9
e/�K���tn�Ω>�818	J����D���v*��?T�
���
��=��V��I��ۏ�_���"���N?&R�ɥjj�+oh�H��/%�{ko��eH�a �@Z���S�	��� m�|�K����ચ?t�U�Wz!6\�I���n6������m@� ��3�~���@�]��} �,2J�/�Q�CklsV/:�O���#�M��j�A!R�(�b�긄.�+�����4��AٌA�g�T�:�.��/��:�~;��{cNmX�F����L'�1���d��|�_���o������2�d�L���0Q�<ʮqqV�c��,8*y�%O	BF37�T��M_x�f*b�4��t҂X�(�����(h�R����;g�ޯ�;��q���g?��@ޔ9R֪^5t3�l �~!&U������HW ���AF�bQ�v.�������ט˻��E�n-xPL��A�j-c��R_
�)H"D�t�XW�@>g�J'_ ���nv�%�yj��2_�bm�L�x��Y�3��^'u<bK��yMvR�!�6�%2��7*���̺=�0�0@�fe�3ďIZǭf�h+t�`gz��X6�E/�ʁNɠe3�-qP�l*����MQ��ӡ)!\��*�����췠�:�O �(7�'`ߏ���\��"5<U����?'=�.N��@�DL+�����"�a���iR�+|�B37�\U���hs@Հ�K����/Z[���`����'�~���c�΃����nӳ
�`�.�1�gT�X�`��p�ǐD���s��I�M�rHD��b^O�a.=kF@�LV���"�wx]����B��wѬO��9�po�N>�ӥ���0h���mUW�2�|���������'߄b~��
RΝ1�?hw��8��߭�acB�D�Ҋ���/�;p�@����\��`��(��07��Y_�b�p�N�q�I��2�V�����0�s:�N$OҠ��`��X~9�o7�A5C%�:�8��]Ed6������s��O+�Y#�����!��^��F��-�S��ķ2�����ͫ<BJn$���H��B�&pz�)�d(6��\�w�Dq����'2���[7�ȢF�3�Y���_~R�%�v�s���-�KG	���m+f�m|}UH����b��[e{%T�u��|ٱ�`�(f��0@�����?���D�V���@�vF��2��ѕ�;v��Xw�޶R ��iުnJ:���F}���\̸=a!�����C�<ҭc�FLʘ���c�1;\4�yjT��r��-� Ϡ�v����7x1U�.G�C;�S��\W)��H��5�:�N��W���
su��G�-�k��Z�9w�[i͡_��y��c����3Y�N��.�%�r��c%���L�I�Me�6P����}��g-jX�t�����m݃^5Q����3J��n����2X)1�t	��r������ј8c��v�޹��l[��h�$����d�����Y[��Ez}��h�ͳ��E���#�s��������r�"�r}n:���!1�m�X����Ǻ��M�ܛ�$_s���"����):������s���wj�=E_��τ_W[�����Bn���� >��t͹=-�ř��~Y �*9Җ)I���?��v���cƶi��E��{�N6�PC��Gi�n�/}��|���w}W�z�g�� �����Ty,�����=�`]\YьE�#���׭����!�tv�uZlT��������ü!�����?� yT�
)vk��}�g� 6���ξRP�||���5�I�e����}zGV��	�ah_�
�J	 ���Z(��ϥ��6FF�ҫ��v�����mW�2���t�t�Y�x4�����%�L��+�a���ٶ�������e�ġb|��w��b�mw�k�{��	tXg�&��d��{g?R7@��g��o�|?<�ξ7����G�&���3woע�,m�s�e�2�?��r#�6�f����$&�[@�P�皤���'�V�X'w�d��*d��f��C�4�j8������:���=�@R=a�����6��������늘��j4���$ �o�֐���S`��ܴu�P0� Sܵ�r�C�x�j�1n͖Ķ[��8p���3s�Bqs$Z�7�ڋ���S�%��Q�i�,糏��7W�qo2��o��S�s����pt��U��#�6�ҡ�����e~�o�ۓZԋ�+��J�� ���zI��Ï��Y��ڰq^ЍQ۲u3�qy�(��cxW� `�.�c�v �w��Ѭ��9|��&ױt��1�[��k���V6{db�I"T�1��^�5����.��Ʋp�/W7��g����������{AQ.��0�Wх����J��[�9p��Oւ@^r
��{K�tN��u�d�����tJGc6��N�G����"L������s�)�0�����2X�+��Q�]����̅�(���!����أ4N[R�����H�	M�c��T
o� �l����z^���\���%+͘۸;Q��{d٘m ^����|��.l�c�syX���Z�m�Р7�v:_مݩ����Y��O�-�rSm��3�� ��s|��X+����4��5�Z[^�س��.CC'��a[9_Tę�'�ݣ& �.%���6�S.��+N�����BC*1-;����1�5�����<M[�2�pzk�h��\ܪ���/����k٪���AzJ�J������+J��4􀤽��¼�E	M��o��˺xa>��/�Nc��u�:{S������t@�{�xr��km��6�ר�{����� �ִ��D0��Z���i�ؓG�8pe=�B�}�@~i)w[����Fi�Z !�i@0�񰼘�`�x�)<�w&~5�ٸuvw��\0�~}���>�ǔ/���(cz�9Kj�ƫ��<#Β�2������w�83�	�oLI���K|�UR��K�5�řG�^:�+07/U!�Ok�� @4��!p���y۶�U=��iM������o�1���9��4Eu��k��s�x���=��|�����S�l��[�PO��7�+�4�By��].)~xn2T�g��ғ���������IZ����iQU)e�T��n���][cv��wxLx�+?}9b��8�篳��o�V���26�����l�DFP���#��lt�������V�7Y9���|M5���B�̎�9�P�yq�:�HZLF�=�@��G�����J��29c���č4F�&{/��Wj؁�����R�6�7O#�y���#x:��$"���y!������j:9
a,�#	�'<�4հtӧ���Cʽ����t+�t-I�]^?Mx-��������1z��@�dP���[y0 �STm���z�����̌%�b��jƳ�n��^��������)�'`/�чO�(7xӯ�?�Z+��v[8��u/�l2�G��Ύ)@�-⮾n����`�;y� �+��{�lވ��v��|��LN��|'YG��Bv�lC�Lۥe���+�r�	��"����g�(�q#�߭3R�����GN�3ǈE�l�-�`�n&�K`�b���K<�b�� ��<	��3z�}�ޫ���d;y�K��!0IC1��W�Q�·,J��iY��a��fo}�|y�?4�x�C��?�S>�'%����M51���g�uG_��7�����.�N���^�7��M?����@�ڝ�K�Q��C9;P|�?,������6�[ߵ���1���s� �:���?��Zӛ��\���U5���eO���d�8GR�v�P_�T-cGΝ��z[-5½1M�^�4��ϊJ h{b��G��
OӾ�K��t+�T1y��sھ�^Q��dءg3���o���������t6"� ��ƅт3��:-Ě���x�c�9Q(k{���?5�3�f��4��3z�o��4�����E�*g��Jc��SM�I���.�E����M
��/�&۬�{�O���-F�]�i��J��᠞ǠDD�?���	p�7؞d�}���?����p:I��ڬ��)K0� #��R��B�#{l3a�gK�Q�((�Ͷ� ��p g�]�)�c�孶%��C��m���E�o�K2��8ڜ�j�<#�[+�U�g�Bd���K!�#kڲ?����J��?���qh�R�<[�Y�X�'� ��^�o��an��W��iI�O�)���v4H�Fm�"U�1���XQ�g�i�[}�R"g&�v&�&yF�
+B��5�q�N��z�2Q��&�6�j�!X�b�#��>Z��:I/�Ą���a��$Gt��$���=�b~���W�ѓ�Km�\�{Ȩ�/#%Au�N�#����,��F�N������P�7|7�v��[ �֚%1~�tg��A��e�rb�������ߎ@��O]MkD�{�"g�M'��7�WtnU���b������$-���-���{
tY@	����Iĩ
��)�a!l���Pw����Md����_4�o��κS�"��̄��-E�N �6�H(�dvP�F[�7�I&ڛ>�kZ'�͡��!F˞�~�	����
��&¤;�����9�[��X�*�z޾q�$ꄔc�p�OZ�t�I�ٖ#@�q�z|M��E]�ifܬ����2O����]� �'$ Xk��� ��%1*��P:��m.��V_Ys[���5�����uM�Ե/ȌJ^=C�BW���He�WIK�����_�l0BҪ��a���,i�\�J��F�j��4[e�S�.�3��Zf%���96k���q��8�H��uk���׼��+�� ���ZE(2vV�(0j�{�)�A�T��HMG��<����l��Ou���V"�����[��G�9	��|��2��(���>�|;+���`�f�˴� ��T�˺ȌT�2�Y��A���EL�h4&�H�������1eU�֬�����uժ��P��Ѥ�J�!A�tT����D��rʬr�st��C�����}Q<|��/�s�X�x� ��4M��G3^Ę�`{��^���ln�'Gϋ��Mܙٖ�,P��b��=U#q�P�r`�M�]�1��v\ U9�@V�~�B%�ǻ���HY����A<OyU#�JU�AN��%ʴ�${���x��6��bq;����	Zs�#��3�	v|8����P����*��|�Rut�7�`:����u�@\j�A��/i��u�;���:e0G3�rl�^?�ж~U6��6$�zj b��a�I�K����%5�.�x��y]`���Vn�9�&�Sw�y2����z��K���Ro�0���8>��^'0�,oC:��6�;����ׄ �J_!�q)K���V?:�6�������/Ǭ1+h ^a]2�x�j����޽���lz��u�-�'`ymL~[!N�ʫ�m.GS��l�JlD�h��>N�h�IYŞ_��=2�nCi�t�p��ݛW�M��P=9?�+y�hL�&b�/����6F�4F�+5�â�t��1)z��c����Kiާ��[�������L^����ӏ	���I�{�a(G����ɷ}��ӝ�Nߔ��nl�3�[ڽnM�L���%�O��d�oݠ���[.�{�4 p',�|��RHF'�]t�P-Ac�����N�V�˰��`F&����G���Mu�AG������N�%%����\ؽ� 0*�#�1{fWA6q��t��K����Rh=����v��-�k�L�,0�џ]��U;��\�N��#Rd�xOv�"�\�G�swᾢ��h}�n�1�f���3����ń�:��E �]����Q4�z���\d�y�~'���X�z�&0뉁<���Ʉ��9��\�����tV]R.�§76\�v��RV5G���i��.��$�BmDiΜ���u�Z<��Y~X�� G��1��d2`6�THv�'���n�<1�\n>�W{�T�� �fW��z��꜄�V2��Y��k����-2*t|И��9�@�]�������Ȧ��<��������ƀ�O�.'r���X��A}��۵����'�g�	^�ps�G���E��T�4#��D�|Y��*���Zw�5�VU���w�2��v�kZI�)w`�]Z�����L�n�*���q�{�I��׷D ���f7��V�-��@?��=�H�*��QY�S��4�k�gMU���=��@ܙ�V��?�PO�Z����8�d���,*C'R���L�1<T9�D	1�dM���1W����Q�y���O�+�f��O2#�U��c��a\�Eυ\6@<�����1��f9}?��%�YJ�,�݀��۞�́��-��Q���4<���RTw�Bn(�c���گ����C��%<ɬȚcc^�*Y�N��%I3��]�&�h�@�W'�+���C%A`���|�|h(>��ܾc}��T��/u��7�̀��.�vus9:Вs{ �IN��Qp�T�rى.���ˆz�f���N?�-���dYme3ۙ�D����p���p:�g�j�Sƀ��,���ه_9��We�k��K���r����*�"�k�ΛH�3, r�f&f�WL��Y�ti���y�Gg&	v�@ny�=�i��A�d2�.�hj�峨A��͡�؉�?]�zvNm�܌�We&�r�SJ�I	sTJPV�YS� �K����Y�ܽ��-s_Jj�P��n�G[��8_8o����y��N�`eF��Q3�ؐj�$���?��16�l�劳���/���!5L�ש�y-xKq�=]� �'�a�!�e���ׂ�f��lsn��r�2	u������2��	=�\�c�)���{_ºO�6�)^ڋ�9> �4�]Q��E��;�!N��D�Z�@��-��wy��UM? n�y�3Xu��!g{���d`���V
L�H�_��`X�߿��W��s��+�"B�X����;ii��,�ו'Sb��d7��W��4�.���ՉR��,�T�)+3�L��ܒn��'l���|��t��?t�V�����K3vbA�����p�7�����YP�B<��PܱX���R[�m��O�;�+���GG��,ﻰ��]�Fky�q��&�ȇj��L�/����տ�;�)հ�����$�B�����X��7b^��@H�\�FP��ro��0F}�7�B6�������ߋ#y���&[/�C���𙐣����3���H��� B�WmV�)8�P�����VI��Rx����75���G$�R��JƩE`��ݜ�ghC}f�S,�/`NAJ9��Vº?������Dј,����E�I#�1Bu�ta/b3���)��������X .�j�� �|~;@�u���&K�u�[_Mk�nfٵ��?'[�� `o�H�,c����f���qc/7�4���_3s���У`�n���멖T��`a���݊`ѩ���"�ܯ��.��9��;m+ʡps=#:H���,u���������$)d,S���� ���B�7��!b&3��5}Q A���h�&��đMsT?��I(�⯫���L��,!X����hʻ���m��Ug����5�ɨ�# �>S� Fo�ҽ^˳�Y�la�M����o�T�dy�)ocM�"Ur��؜���TCz\�,���\����߹1��I������;7(!������2�߹�����܈���wn���������_u�l�0�/T��uҰן �� !�^kK�X ܁e[�Hxǡ���I2~���5M���8�@A�8d��eG8���{��W^c�N�j�tR�z�u ͎�@�<8 
oTd˖[U���{Wn[C�;���$�g�Ʈ �&Or��<�������=���h��s���T��%U�ƜGi5�i|8�?�.�@'�!1�XY�q�(����hX���+�iR��l�0"J�	��<�uT��^�'ԝn�j*�9���2��#y��a�D]�q���Y#|�<�4�$P�d'�mB��|��i6g��A��������Jɀ����|Xyq�f-oBK�j��)C���ąo��Y#�@����˝Ҕ>�]a��� w�tF��O_f��{I��`;������>1���FVH|r�
EK�-)D��+�䳞��w�VJ��CG�}���寀y�Ѷ���5.:���G7�:?j��_j�����_�A��2�&zpl?	�9�F���N��[?�7bҡLh?����5iPÛP�c���n3�#��16�����	�F�]{^���(�֏}����ւ��`JD�A;sL���N�,����6��sw�eM5E�_�m�}�
WR�1����7����z���u(P����ڣ<�W,.c��)��/UǷSQ�������~:�d�|K��F����6p�m�OE}�(����T������
���`H�h��������L�sS�W��+�>�����\���
��l��0ê>b��M"�b6k�e}��M+ҳ�R'ㅜ��F���^����]���n��f P��B$���o¯�oP�"�@ah/����\=t�z�+/�<p�+)�!��y��zȽ�1nn�N6���`��mOR���o�zT�ۿ��C&K٨-Bp�O|�8�ŧPT���^n��ߒ/�4�T�W|�92���yEV'�0�,�q+�т�l�.53�{).��ܖ�'O���>��JO''�8z"�	�k!D�}�~�~'�s�%}�W�T��ߵwst�^{ጣb�k�,u�$an�!M��.I�-KT�Z��W�Ā*����bw�ն�ȝ�����7�w�i|,�������=�A��㌗�7�l̈z�T���;��������Rb���|�8��=z ℡�	�F(�/��H�ЁE��x�?C�������}�D�M&n��=��(���x1��^�B��I^�G\�3|,ݦj��vVh�M)@,�I�+e�"B���c�)�cmP���8���@�P�B��zlݼ��u�+��5P/b�c1M
��l���>���,�d7Bw��ޏ�:�(HKyBm�iݶ{]`�"�i�1�ftN`�,"!�cK.�Ya/wmm:_N��·^M�Ţ���t.�mo�/�V�R�Xa�xQ��4��<�o`�X��������{�9��+m��{�����Ռ
&�nǢ�VxE`���[����tr,M�����c�DE�J0;%�H2�>�t?�x�R���F�.Г�i���q�܉��D�ק�}RL ^x!��)�8p�<<@v�u�� qG�����4S��@}�t_m���
P-��8�D�@y#ý��W3�K��?�f޵�u����5������s6��@%�-!��%*h\�Y���bS�T{ܽ]��O<�{vk*��!���}��^?*0�Л�p���0�y��ye�`N��3��)s���>��2ݱ��=� � f�?�)]�lҷ9��1���j�a�%p���|�̉�F t��<�$�0��r�`r�奷#�$�x�%|��/���ϊ�@�n+<��l���VB�?v��(�6��{���]o���z�������@���?�UqU��<d��M�P���}�I3�Qoݸ��wgs��'Y���e�.�r�ވ�n~���	6C*,Qx�T��i��	c2y�õ�S��s����5������}p�;XJ���}��$v���'M�iқ�4L��PxrZ��j�^h���?�C��!r\�I9�z������2h/��N��L8vj����.,k���џM��Yv�����VԓO����x�|��5�"�=f۷���KV�M��$���[Ž�$yy��i�*T�W�(3���̫�EyAWi��*1F�Z�+��R�D�Z0��žyl�'�z��L*���ڌ��ٶ�`EV+>u�.
;��������g��g������5ȧ[�
ߎ���56l��(��;���mw#�M_��u�*y9��(��2�?�pP<Co��-<�����"��RZ<���F�Ϣ�"�wY�~i��`x��b������X�\�v��ɒ�6�c���µqh�\��{��b_��i{�硾���|� �6�-�f?�.O^-X�6��:��=ZwTP�������bJ�J����ۚ�m�]_�����{Mp���,Y���jAz��G���5/��t�r�Ӗa*u�N�i^�H�Q�?�$�[���H��oկ�p>���+��vxk�Dё�]����/�q���x�r�)���ڬ�KX�`��G�~��7S=<�1�K��0�E�Z�#Du���Ӿ�\²z?��{�=�sNE�f��>���}��eK�!T�);��}����Y]���`J5��e�B��Zq�z-?ΈO[0Tc��ԑӂ}&�פ���7u�Vz����'�&��;��aR4�������Gqֵ穖��sa�x"m��`��IM���`�:�	3�s`z+P��{��̬��˾e��W}oȫ�΅D��j�7%�^J�鮷$cQ��\��^�$,0���C����N���+���;���7����@�na��dUbqt6���>�����8�y���[�h;!�/���?�u�+�"���g�����a�y���Oɾ=�o,��tV��h[+E��`��u���j�L������R� +侖�O^JXOv���#�>���~(��켆��_������g�}�]���.��g��`s�W*ݬ&�+�t���cZ��+Id��x��ހ�@C�V�E�Z��a�I�%���o�N��)�MR��@��)ijIXV��J�h��~�ΦM�����2�ݮ:��8�/�7K���ܟJ��=�2����[���a	��;�5m��5-��QWj�R��d�O�1
z��DD_�B�.��貸��8}q����&4��}T*���=kj~�q��|�+3W%`�<s���ߜ�T�r�d�'>l_��� 5�gSP�X���u�	�`z��J:4�*���,�T�5m�6m;eu�F���P�8�*d.�ꦠG����K ��D�fmO�lP��r]�&e���]^��	C�l���y�`Q��4����N�M�s��2��S32����k�b�7㖩Z�V�=5����~�ߴ�>����5c�ewc[�6y���D)��,��O!�v�Ijso�ᦸ��Dj1:q�3�d(w��.���W��RX^�ws����on�hvT�}�xG�q�S�ě�C{{J��!ώod�a��D�>��g,#Eݝh��sQ�fj��E��V{�k�N�"hp�A�#JW���2a�ba?�lj�b��R�5h��{�O�oǁAwEFWQ��8��8�_w��'��$�ww��A��;���r���bB���<]oIxi+lv�%}=�e�,ҚN;n�j��_�L�d�"���������U�����+怖���'̸�w;��6#@�\���I�[��5��P�%3$/������w4��s
��
��x�~�h(�͢@՞`�T'���<���pnI ��Pl`'+'�� ���XӶ�[F�֍wفO�|ʠ��+���q؃��%�ٍ]�����̏&a���o1c�ɐ�����T�/��ο�D�d¡�(�3؋��s!w�B�6͘{F��&O<��[Y�w�F<$�ME|�5�ۿ��Q�5M!L��зLL2~��b+i���Z��hR�?�t
�+�{;�w��͎��m��@����/U1G;�'�

ll[^G��?��N_z����±���|aCg��a��j�x�Z��x��n�+��|e#=Q�i^y�k�8M/[Zǆ��6���B<�A��i�7;n�z?�y��������X[��ʡ����_F�lnv���$�i���~,��hw�sN�e�m������۶�allû��"S��f���F�ҧWa̷���X�����r'%�O�����r���|G�Sґ��n����HW,�w��N����i�QI�!�q�u��F��o	�h�'�n���oEu>A��/r蹲`��p��BB��6A'X���m}�����B.���Ħ�eC��W�Er��y~��#��iW
�&| +���ڵ#�gg��;��M���v2�:<�ܳM���4w:ԋ5���g��Ev�����Ք�I�:��m�h*N�:M���D-��E���FW�W'���t�u�/�j�D�=Wc�!�Q�x��%u����E�JBk�"��V��S*@B���I|M��?�0m�5vHn���cM�I�$P�& �9�C��N����*	�[j�%g�yUj8��6a�L?�T\�u7��\���T�'ޖ�h{�r�4)�lZh�*�uu擓�����l���C�}���X�w�9I��ON."���h[Ph�	)��Q�LL�����,���7-| ���9��-�c��?���l�����},$>v��z6�F0s�`p��(���Bt�~	&�U�#-�BS$t�Z���u�#ôɴ��{]�PF�Ta-BO��` �ˑR59̬�Z� � �6+��S�ֈ����tT��[����ޠ�0:�Ԁ�����$w�a������©f�������"I.�T��\����Q�oz�&����{��1���|`��^�1$�u��f�)��<�� /jܳ{�k�U`�D_c�&F/̧�,ȁ����a��k���ڡ�x��o���'Ɛ�C`6���\%���0��6
>I��ܾ�'ro��Ro��	���U�F��jf�&��JC��ow��h�u[W�)G�0ub<�U<������!����ٸɌ|dW��5\S�۲�^(� �(I�P?1=p���'oC��u�C�/�Ƭs��Kk�{��b�`E�;�H�(����s��\�a:�r�[j�!��	��O�� ��s�rd�c�%*dݒ.��8�Z�Rk3���v������1��~�_�_��+U�7
d���2p��?Pt���'��Hwu	�L�3������7A�Gk45��ߞ���=5�$���_�]�!���b5����Fn\��n�0�<r����˹'Le��տ��9��B3���%m<�^ly�,8���om�ʔ.��0��x3vh��r�E"8�yY�/���0��S\�����n�8UM�v�9��~|��M�JT��t�uB���uS�S�IB����������8���~��S�9{�Cͫ�P'��##�]1�
�P1z���x��iiq���񆼠S��D+gR-�Iƈ�qơJ�7��c�O>����}���咥x6*����!��A�b��k�H�F���N�����u��(za�%�>���(�PcñZ��F����^��QJ[?�ZY��)� �y�����^CL�iW��Z2 <x�_�;ip���&˸x�>u��Gp&Ņ!����d�O�mgr�l�VK�yv���E8�:��sV�+cu1�?�{���$���D�9o��v�e���q�פ�񐨵�&�nl����D������+��A���v<���0���Sf�������Y n�'V^J>Ā#�~�N�Mu��<�@��i��s��{���]�*�V4�����E�F�I�y�� ���� (�b"a`H�,���GN�n�
�jcG���ĨbHoV[Qf$��*n�4��r��U>�LJ�m0��P�����S2#C`ڙP`J�r���[m��t�"�x�.1I��`/7˘�Y����
�F��Ep^�lf��Y��������99Z(����2u�e�CI���7�&KSG���HM��|rz�~���(\�w�#6t*�r�����6=�	awv9�0�$x{�#0x�o��>�����M�����I����G��kb��D�oH��eC:�v���(l����E�jf�H�`=����������%���D:7�  HwHww�t�4�H7HK�4Hæ��E����s����wv�5�\�y���\$�%��I�h�7�]�"�Ux�.P�>�wB��ľ�5l�禯���{<�mm�*K@��B�2B%�DBJ��B6ڨ,~j��u�� 1��(&��h 7'�/E�z�o�K�S�#j\D'%��
n��$���]�~�]��$T����Jo7�eޙn-���a�h�L2|{�Mo���K�7y=��o���{��<w����F���)$(���<��}�*U >$��ޣ��M��s�	kk����'�M� �{�����S��V_��c���CaZpZ"��]���#>�@����;�jbrK	�j�cCڿ)���xoF����� �pM��o-����v��Dk� +b��T���X���Ѻ-��s_��Ӗ� �K�����+�����.)Of�\:�.�}/�����8�g��c������0��w��8���L�Q�)f��>��¨��!`�7�6�I_ h3�4Y��CQ3�SZ�Lɏ/m
!�����4��Y��(/l>6	4�+���\&�N�G�����4�q��Z]��Ӎ=�Ў�����-,�ZA<����9y��G��Vo���+v����02�Zv���v	��5�\$��ڼ�a_Wx�>���Ks׷,�ήm����zyzB�B���-�XLG�cߖ���^�4��R��Zj�NM�tj�uK����d�@�C#GlL�s����	 � �Ԟ�f����>���6���a�����h�wu��~P , ���v_+�"ۄ/�\y�_��XH�f���m���M�@ʂ�n_i���%"����H��	�ay	,���g��'u�O�ɍwr�pĶ�W.Uh2�?⃌���WE�e,�;����e��JR����,���nxoP8�p�$s�;�F��44Y�k#:�>ַ-��%��'Vo>
��˭�"by��� �S��������p�Ȅ��sg����F��Iv�'�=��mS18�xG��h�y�W�������eB`�z��D&g7���Z�CQD>�ű��������P��b��qjg]#u���i�����ō��d�"������>^Fk�����D4Oƥ�Ҽt��Y�.v��Ƴ�I�<�B�>חV����Հ��7&��޼95���l���	m^gީ��l&��`;:t��5q���$��@	�����,����M�����_���5��XV� ��'>�޸���}M��??�؞l>R��]#ML��NWf���� 4H��+Y>�������Y�]����ڕ��4�-Mv��X5`�1jր���I���(| ^rܩ�I0���aP�4�+O��Y��geˎ�b|u��|;q}�����!����I�z!q���4�rbo_礊���1t���e�+PKtƼ��:‰s*R�\���ҤM�	�Ep���1f8 �������U��A#��%�{eQ�.ޔ�r��!)��
~}E�w�`nͥ��dt������,�'��k�O��-�MY=���y�y�7t��Xk�P�vpm~:bc���8�����ā�j�1��N���5P�j�]�������w!"�@'�o7��4�_����E�6��E2xE%�7[� ha�|��=^��S=?�ƺ~��Ex(��9#�X���0�m��	������{Е$�~Ǎ�m���+���~Q�W��ހ1(�τ�q�5�t���z�t�� ���ǾlP�Q���7��ڋG�N��xN������V�����o�	�P�흍�{d.�L5p̿����Y���%�t���J
��p�IU�juBC��X��;��׮{��A�9!�0Gޑ]�\P�O�?��4�)sG��~f�!R������X�o�8�(Q�g�Ƶ��-�	F'�z_���G.��T�Q5'������A��sC������3�H^��+[�Z�;��DˬP%:�W{8N�h��m��� ���½�%e�:�OhaJ+���[��j����.a�"H������:2���6�l���� 	��6�k�sQk�Q�++��{*�{���G<��N���o�̂e{yW7@4r��Q��P�-C=�OW^-�f(��W�%��f����K؆��z<K�M���L�s{=ن� '���7�SE&�w�����������L���]M��@�����,�%fB����<�/R��$t��b�kQӨX X���渞��u}NG�	le��+������/�ǋg�I^�+]�{�A#a믲x�׿��:1��,Q�=Ձ�tCK*(b��s�w~��Ý�w�k�o�R�7*�/��\!�1�ݸH�d�^�VS�=v�m��j9���C�RE�Oϩ�w�K?p���"�]{B��HHO��J�.���o,�o'�͟���ӣY�?�f8��`d�x*�b�3��*JAr�_h�a
!�Ft ������)��\Jz����/"� ��D�7��z��2��*Ʃ�"�����KV/�s��(}�6��9Ԩ�r8�CԵ�^��8y�?v���(��W4�1Cl�R���W�U�.��)ó
_=;�z�5u��&M�ߚY6C[�2#����У�#?,���#�5(��H4��?��l���c4o��B���ǎ�R6�4�h2KJ��K�3'�:�r�LZFG�f�5�1Y��]:�-g=�%��3O!>���`:)8��[�N*��S�rc�$MVg^Wm$���C�mf��1��,�e��A���a�
X�-ѫm��^�Aa��eQ�a��k��( ��ݜ���dd��P[�j�bþ�y��m��
_��z ��������*�yQ�(�d���w�M���t,��Qk���e�B��7%��M�K����'�xȯ���;5�����+�m����FCѡ�ߓ������������w�pފ�F�%&	��C�O��.xە��o�O�	}@��f�%�hU:�pc���=o2�!ܛ{���!ʷ�"���w.ho�=KkO�|�|&����ݭ@r������ux���hF���x��V�'C���������Z�}L�=4-ʑǺ���Ĉ�ţ�lZ�,<�y���E/��6��ߓk�v�O:V��]������E���w�Ɗ��f'�*B��q�����AA��������N�$R]��W�H-�4K���� 4.:���5s�iu�#�}d�[@	
wv�s���^�u�_�4�T�L��L��Q���p��;j��*O�U;����͢NU�ӕ���c;�w�'�Ӫ����H��F�L�:Y�;3VC�l1�S�3��	"p��s��]mտ�����n�9�(A����K�8b��U%�@M �:��<RV�ni.����z�xGڥj^�P�I����S��3��~�����I��asFX�V��~��	&|Y�p;%��=%��,�14��,�9����=�K��%��ݏy�~�]n7mF�Աσ3�R�)󎀤]��q�e	��io�|���R7�?���x��e�W��(<�.��Smģz�E �q�׳��/@�˳b�
�`�N��b���Q)�Ӹq�35�;2��%.ⴰ�KGw6��[���i�Yɻ�,����5
�7��������	�J�h\ 
���
��~|qWgLS=%��aGpޔ�H}�<��`�Pa�u����� ΀�%�M�� Q���W<��˨�*�.K%K�;��3��ǫ
�^%h����lEy%6��������c�m�-�-��|��2���=�(e��bze� Uh"�ɸ��`����9l�0�\og1g_�
V�Q���ƫ�
?�x<�sk�������>Bo�\��A};J���&�%d��a ���o�ZJ��̐|3`���_��t�`�]�~����7e��ҵ��g�.�̇��'o�� �����́p>*�$H�0no�F1���(�!�Lq��|�YN��Fsg�����2ٲ��+��$eJ�%�_gߥ"Q��A���\�n�u�"�?�L�z�T،;Пg?�8d'(0�q�\g�3��>��p�tS���\�Zr���B��d'��>~�X7��5�����e�Ƴ|UOO��f�/,��M[`����S��̡���g3QS������'����T�@3�L�<F�*�}'<����5Z���y�=��K�w>�E�$q@Nն$e�^��y��B[�M_i/ᣒ<3�Rk���l{�3^���L�q�NS3 ����v�^�{U��D_�����Iy��@_�p~���ql8��E%�.���g����ī�n@�d�'{�iou��5(}�Ӳ�qQ�
�j���'�W�'���1���M/�x[o=vL)�T8����er%/�|G� Df���;�,�&k�%k�o�ɭ�,<��&���K9����;��Рs�����D��T���R���U��B�(���>i���(��'S�l�Y~F�զA�hZ��So�k�&����ˋ���M��*�� É���,h���d�ڰ������GuJ�.?�eb3*��mo��(YZN�����v&2Q��c,��j��>\���;�%�h��J�ׇ<�������y�������tlD�'[�v��6q� ��(R������[�qa�h�m=8*�����f�fi�N�i��0o�]#HH�仃���'�/�~���f�h��;��S����c�m_ݺPb�oM-�����#e��D��p�M��ֽu�>m̫	�3l�}?;�w*����v>, ������m
�#TӲwkX��M�u�i/��!�׈io!T�D ^8��S�sP�V�q��i�]�xFܬ�D�~��Ԟ�tjR|���B��b 0������(yq�e;�T� ���i<v�����4�3z$zʋ�[�������J6��Da�	$m-PV��i���Vn�ܧ���' �D[Tfw�e��{���m�H��v��-Iv��2&�����VJ!nZD�����A�xP�c1��,�^*lu�����s�U�F�p?��N"��?\r���jG�^��A�=���ǞeV�8�5�\F �U���{ݚ9�m��ԓg��"�6_�bpR��w�ߐ�J /C�_R�1�Y��j���-��zݗ�pA�*
s�Z�y�-l	�.�Y�U���iLȃLr_�y�z�w�����+>���R-��̝�)Q,Y`O�#��aج���}��+C�W,�	gvK{�L��]c��y�c$o�BGP ���I�ruo��`���MI�a;��s�ʩ�v˥[]`NwDP�Й���}MfH����8�\���n��"aV�+�ح��S�������qt�	�^��I��sH)~�\8��Һ��`��:���u�a���)`�j��eV.�p�w�D�T`��w-Jfv�N���=}h#Kn�Y�W ��N����L�ߓ�N�9\�=B��d���B�z�Txxh(!̑'78=/˸;���<fW�v�-gg-���wz����y-͡�f	�n��"V:��R5\��F��F�M����\,_ݖ���ܽI�S)���;��U�?oaI;�8�ZB�&M�C���Ж��5:Ya������9E�Հm�66]�\`�y�w<H�+5P���h	@�a�Z��9����y�����|�K��[3���ډ�b��A��Z�X��+�ǩ�׾��kL�L�T�TkGB���j8
�
�6~���G�����p����M�d�/�h±����!�����St�jp�Q@��B���ͦ�e�d�&��&̳�
�Ύ��I��.���~5{�=�bj`"U�S�g����Bd`Ok���	@g;��W=j�!^P�Ӆ��zJ>zA*�s�� K0ֿ� �*������Xn`���;�b Z׉c{�ĸ@�4z��<���c�E��-�J{�(CǠ��+�F��\=?�2�+u�!�	#�VO�(�	L�tNf��q�r�z�	�=�<+���6�~� ���~@�8A2��;]c��x�@T�;��Vn���Ը���K�20nt 
Fn����ElN��6@����L� ����/��]�(�!⍱1��O�����{��V���da����%��"�����Q @!ʿ������|��t��ovD����~����V�g�X�+��B�\����<�t�vK�mq�m���[�rVn�����	.�`9x�������{��:�+�t�,*L��/o��;��`��)�������!|��HF������h�HO�Nƨ i=�97����nwڸ��leGMv�ۊ,Z�f��#CjE���.|먓\H���@���߉[��i��ks1A�TZ%P�����'y۫>�v�^���_2v;�ة	���]���6��⤥=�|Cc�7:m�\��~�#�m*��CJ��>���}iI� j�Ga`;^�?�%�L��D`�W1�wƁ�%�DH|��vަ� Z�@,�HB=�����3�����w��Qh���1w7n�gN�C���s�c�z�n��Ф��]��H�}}�o���⿜�� �3��,��)cL:���_�Z�V���]!	�����C�.#��l��p����v�ү9I�ؓC�F�_E;ʍ_�툈�~OdH�p	�*�"2)	Kg�/����&~�[h�̠K�A���m��_H�]�s��`�;.<vs�&�7�^�g�L�qȕ��	;�-�<'A�{��緜�u����0U�Q@_���R�;�az��c4X}�:��Ii���j""*��.ˈp�[ߍӈ?hԐC�W���Y�Z6r��}^�b�����V]�Wo��l��D���=Mځ_ӥF��'dmN��7%���E���7����L&"�~�ژ��}��瓉d� ���m����fK�9�<pߕ��*<K/��M 5Y�4A�����%��	���d���s��?�6$)ޮ��3�-�)/2�{�荐KxZ��~8�Y���!x:l�8!3.ی^�<�5�'^�W	M��+S&�ѡ���Y�@M���M�Vj���w�'��<�i�4���oq��Z�ԑ�z�4�L�a�ϖ����W;�d�۱B{�Aap~F��(��1�"�o�kΆ�X
Ӟ��\PW�y����2���4̿�
"1�ʔ� Dl��&��&��
�w�h-�ur�(_8P6Xj3�l���D����(�d-=�C�((B{��PB*���-M� k��M>��a������ǡ��Dl�d/�0�������m�qt?8�pȏ�.9�Ҡ���[r�aptc���󺡡������n"��EBW]�)�X�ge2>@�6�^`���Qo�o8^����Sq8d�vIӣ?���޴��"*صG8��-o�����ʬj#ЃP���*�l
��(F�k�5�S% ?�p�郌/8�Q��I����+��� �N��m�ݤ��4�ى`�ӈL��ڡ�I��H(��k��Y�0����	�Tu�Xd��,��ڿi@����w��ی��/�͑K��z��Y��F?������J-��_�T��[�%�z�0��V<B�\B�ȩ��o�%��Wlg�����c���$!���%Pi2Ns�  �b��dsXA���|�h�U�i ҮX�Ww���
�o�Bj���s���56K]/�վ~^i$?���S���d��7ʶ�Ksj�r���.�L��2F�7�	�P�z�f)��<���S�Nw��ڔܐ��\��_=W������Z�Ƽ���:�b����]B�YD�w��qP������2�>I
ă[wjEuv��휱2��Cr8�RI��G��� A���o9��ԄL�&=n٧3ZSǎ+ec� ��97;���L	��5��7U�5���2Su�c+�i�dg��xT?6��QU%�Hz����8|;��\ւ���\V�hJ>��'��$�-v��d� �NtMR�m�l,		N�����D�a��R<%��M&���*���c��9�ENz2�c�JD8X�]�G\�ޝ����X�L}kbH����&�ϝP}+-��yhJ���u::�
~
���Ú jf��6�e�@�EN����A�cS�Q�8�ߦ���d���14Tk���ݺ��%�Qt%X6v�M-^�YC���$Fx�H�DH�|N��[~����"|+1^�}2��2aJ��`/p˱�vr��>���(3�&���G�m�0]��l�s(�䰢�R���)�qq��J
Gj��љ?!�^X�7R�k-�⹳�ԵS��$��#ލ��|�%";y�����������?�׿�g�\����Qw7�ڪ�e�����硅��5���^f�~��ً��GI������.c�R��G�㻇C��d��%���][RH����
a_�$�;)Q�v�]u��{����ONWww��P�����L*'h:��@���kV�ܞ[^�������jZ�y0L8�bş?���t�k�uh��!v�F\�oڭ7@C�FHJ7�6Oj�U��9@�;��K�gw�b�o�#3�s��rv��B"�./R�d�'��m��T�qE%�����n��J��k3d����:���7�|8m�|�?4�L}|;v�yW�bq��1�v���ţ����A���W��"�L��xJ�h��^��{=L
�o==<	c�����\�-���n��-���z�-*H�6[�~��e������Ei�F��0����՚1�����*ע�x&���/�,I��b��K�$�v��g�I.m���g���^�x
���S�Jî;��@$��lݴIzJ��O{�o�ʾ)�S�j���K�K�eǁ���ʓ��T-�>8�;���w�jZX����:���S��'��R=��ے��l"v ����kG��� �n��>����u�feH���g�H�O{z��2R��8L��ct����GL�V ��S�u��7��n3���X^M���e�"����E[���\�/"�ɯ���8�U	J�ܬ�r��D�F����_Tm/N��'�N��0����a��K����1Y���*U�eEG�f����T���^��'GP`�;x!�\��ق�Ηa҄ E�"U��j���X�O]�x��$[�(y�Y�VQ�p�G[��F�2�&���D8��0�/"�˸ 't[���	a��A�pO��'B��!$P`2/�/���/ڸ~�m�rO�������?S�9�YA���w��2D}�]E�Ǟ�N�/�`��P���߈��יƉf���o�Zn�����[���C1�;Ǵ4;�w�5'|�x��0�	�q��t�אZ=}Q�d�O޲+J ��J�Yt������K��{89�<x�#{��Bb3�ޟV}�B`OQB�L�:!J�<p����q�*���yP禿�����㊈���,ٟ�����,�9�t`{J)��J�6s�R�a������,t'����XX?T�������Sa=Œ��|��O*���r�Kڃ��L�s��$L���8�s���n���ξ�h���{�K�� ��܄=���y�z�|�z�Ք�p"|f���D6��(ͫ�q����k}����4����bu���~-�]����0�J�95ԄF}1�D���#q��W�~1�jl��l[!*ʟbӢ	��=?� %�[�����M��V���Wb�w����%��n/v�J.��*ʹ��BW��Kpߡn젡�L���S�nD�A��CV ��r}C$?��+EEvR�s�zr������u¿��	�i�̲&xU��o���L���:*�OQ%�d���U�h	=���s��A`߾>;���.eʱS�0�k�Lߪ>[2�z���"� 
�f}�����,?���ɴ?��0qLih��x��#mP�T��ߋi-�/H�K O�>��2�M��X�wmI��<���x��V�y�Ew?ʹD���	���T�l���<�銺�C�osG�^�I�Uxrl��\�4;7Qw�F��b��#�VEFfm�;q`�J�}G�6�c�O- OD�0�k�Z���8�gj��D�gHk�Rڏ#ΤK�:���W��~�m�\�S��2\�%�
��.���S�؜����0It&�������G�d��U�ҋ�9 �']�������o�"���;�cC���j4H-���������S�̵��c;v�H���ٳ�t^	��T��g������'V�	{����RT���GB�]��ؘˁ)9�b���E��-���,���ɷپ�Q�$���b�}L&[~�f�q��ůY�z�]O����X�K2Κ��R"͞s9�����n�h���{J��k�4��	��a���3��(?���?��6w-5�s?`��}(��n����;b�}���a�#��^z�XC��#��e�ϫ;Z��;4Y�nZ����MoH��֮ݭ��
-�EmW(Dn*Q?�<�j ����L�]dހ$rz���T����h)ϋU��1��K������h�.x��~�d���Ĵ&�*��x*�� ]����X� ��|��_ɶ�3�yxv'�byV�aI1���8������n�|gm����x��N��BsϠ�}�٧ �7�ς���'�D�����y�����|�7��	ۿ<��0��>�^	��<����;�R�,U���O�\[yvdaJ�6P������)��jL�G1�o(b�.��+�6��AY._uS B7��ċOfs�E�Wp��E��=�-IEKJ�hAe޻�1�OYH���@��bJ�t��S�c�U��DiC{�`5ЄW����>sěT*�9$��o�J���P�rdj���(˸{L$�A=ޔ;ȳ5���;��@ʯl>R���R�~��v� ضϟlzY)|}��peM?�g�5l�H8C=�R��3o!?�3��/LH*+
� ©C�w��n��IF�S�/;�\���w)�5�T����?��?t���s8$"m�D#�ea:��p���(F�O-�8���"K%�;�x̘�h���� �X���R�=p�T�W��s%�Q�9wm��7�L&
c�'7�4���>���r��Z1�����2�y���X��.���+|?j�"�\��έ���d8�&}��})��``�^$�5<FjKوs�w�����ˋ�r�ͦ[0�<^{��-�OZ}�gdy���x����0JQ+:Gt&D��, �n�ݾL�lz��}�b�0�9�C����J��{qlkY���]��XvW̩�޾E�\�쑧~��Vw��Q��P�b�� g�q�/��!��	XĈ��?�O#l��,7i���_�\ ��0���Q�h��;���hZg�e��$��6��]�Z@z��f�i�Ov�M9�7B���%��js�Z�o��n|�>���c��~ӯ�:i2f1��'C�ܜ%$����%�z\�EC��~Cᰁc5�������X<Y퍔�(��Ҡ�p�I�=�ו:b����	����E<�#��[�-�p�3>�Sw;Rg��*���u�"u[HK$�A�����oF`+S�1~�ʢ@*��2Ka���j�L)�2�Ct�*'nPM|��X�H�����V�/b��$�6���Ǝ�!P���J��h�i$��͢��H)`�a���a�_�Z֑��.I �C������Ú��mdlrJ��:�z���94�m��������Aȩ����gă��v�ϋ�N�i�j�D:S" ���*��P�ң1�30�cO��Dr���U�#��t6k(Rubd�r}�ĸ�v��17�a�
5]~��$��c�74��}�y.�eݑ�}����A�G,V�+���et?#�뗤��֓&� ���>+a'b��6�P�>�lc[�*�W;��[@N4`��?���� �2Q�ݗ�_�9�R(Ͱ=�Ő�V����_�o�)��J��	�o���h&gn!����=������6gkV��1W14��^Ox�(O湺�C\��7��k���f�����̩Ek�+�@Ye��1�F��	�+��G1D�@��0�!�K��[���;������}�F@Zl����Y+������e��]���l�q�6K�f��,R��v��*���E)
�e��:�ܙ�ά?_h!�\-D%�HZ���?o��� �	���,/��AT��EF��D=�:��T���,�z6~��RxưE�P����e6�kNKɇ�[.2�{n��\���噌��sj6-�������]3O6�E]�ų��T���,��a�|i����ИMQ����ןdɔ����Q�MR����l/?[��r��E�����ȑ���cL=��*�`fɳ2���۬Q&/����O5dqE��}��m��=���5	H�����l~�x�)��):�q���0��~G˱釻����A�'����|H�>�U�Q׉+/-$ ����^�%؋y9[�׃�z-�5��R�����p �gix*� ���m�Z��
���nӥ�Ryb;�Q[��F@q�5l���~�ō��UH�nw�����~5���4��-��^UJ}�Vx;U����s'�oT'��Q���b}D��!�@���^�X�9�c����uQ����!姊���h�������j���k�c\�7�N�G%�.�O	+���|���bg���k�F����3���\5O��=�协_g�V����h����[��-�0b�9`�i�S}w��{w䈿.D�*�	l&�|�2�P������h�w��7��&'$طN�ڰ�ն;���w�1(�󔎩sI�\�PO�f�G4lrDgAZ�!���o2�<�;7{���ݮc/iGU�޻Ė�=�r���բ�/�ۺH:wJ���	P�h�sk�� e��:Fg���	����+�� J҅�e8���i������������ 8�U
1K75��Gt��Oi��K8����^�cR&�K��)�mI��py��#ꗫ[�*�H�y����f\�����Fl{��2|�i- �$@�]T��^�/�d]F��gޡ�h�~_9I�ǥ�����~� �߾kY�i�jȖ�-^rD��T,��#A�E{��/JC��}4%:�©�w�ϡȐ��5�Q��|;[g�6d|������>���c���k���6�.a�j���+o�
g)vғi2x0.i_��09����iM���·㚩�*;�ܞ��{���"'>FA���ߣ-~��櫦��OC����q2��}�B����4�f˭}~�Wvi2e���l8H-����Iu�=�� �W8��p�M˸4K�x��vH�pY�����ޘ�oAJ'J6��*����)��!��W!���KԲ[޶��e�[p+��o���A:�줪�-�;��HO������&�I�s�{��ubZ��/�
WcP\�v
a��#)�?���X-���^�-����F�'y�O���{#��8*�l��PA:�v_6��>�r�l̬5��g=����jk�@����W	�7�
��~�")x͂���pڭ8�BM0\3j�� N!�E�H�Z��L�������p�tɷ��*�7�	�.��)���ƒ'�}���!(r��2.��E[`�h�*H4ʬտT��z�Й������v��P�B˯��t��t��d!�G,0*M
���ܐs��{�fEkίc��Y5(���ȣ�zﾭP�$Slr��"&�9w��҃i��A�~���>�6���Q|�tƚ ñL��V$�0ZGriy9zL����z�l?��X�*��H�?�&���LE�3��]\k�b�(���e[/�����4�O� d3	!��d}��[�"=~�ʳr�c�1��=��\]��Yo�fō����~��	�NAAj�"�VǫV9�����>c�\?V4q5��u�q�\��y:�>\i�;6a!c��K���������Cha�R�K�Μ��
5��)�Rovvz�emj#��)x����U|�i�ʖ6��od 0h���L�4c=4��i[�w)(_]..5r�H�/�a��p���\Ѯ�HU�I?���&.>�$�a(��
@0����C����	�?���*�������w��}�����G����}` �
�G
_O2���&���#��N����I�Y�u~��������q7������o��R9��Zr\>��=1��ds��
uw��n��U�$�s��v���:M����NS
���D6����4����:M�@���N�}���,�����4q{B��������K��_JxL�����`�l((���겪r	�6"���əި�6�w��t��2[�V;q��p��<Kh9X?wP�Z^"�l���Vۼ�O��s���U���a��e��	[��gde3�5OA���ZK������������"��Z�y�-뷝d��I�z�
	��r�R4@е���\mas��?d/֕F��ow^�|�uU�0z�wc�����gI�X�V�l��f�A#�=�)1V�h]�v�D4�CN#>22�����7�{�!��[ג�ת�*	Q]�Gq<3�v{��^�D[{~��ީD������\��K�6�u���$��r^�r��x��?�O��w	��>�Jm��屣Z�L,Z37F�@�9b���(,Y�~L�)������+r��m󒠼e��UVp��j����>x�\��T����i��ɍIH�/��AC�сZ_W�~��dC�r�.+�?o2�j�Y���a�S:N��Vv�
����4�����N?�0y=0�u֚�$[|e���(H����������kIs�2}5�
|iBx��"zyڏ�B'��e�d��a�jw�{���UF���߂�����{4O.����7o�,���?T�4�"�C�ߑ��Ȧx�i�q��/�>���e��H�1�YK���4�j��0�H�*�k��
?�1-�棼�"UeI���
W�paӹ�'x��p�Ǣ�0��և��_�~�J}Q'�x*8�������8��v��m~'y�3!R��G�v����7���(�[[���g��\UJ�o����H.�Hh�t�ֻ4�:L����?I�P���Y���.(`���R����f�
/?{v�K��%��Dl�>�xG.%�n|�#*�I�g�7l��Y�h1vE��Q���p3B�:����f$����k`�$������}�3�\|��]���k�B?�z�&�7Bj�si�¯�u7Bv(0>nM��Ʀ��5��%��߃$��o�����#��e!yF\ߖ7��cћ��?��9O`�����,�,[g~+E�����)����H�p�K�hՍ6��&��h?��|e.�b|�-ɿ��0����D���k��v�����~*���q�� R-x&b�GAX<�B�A��������BB����O��j�a���v��tg�w@Z�Z¥F,�1)��G�Jg��g�Ļ��KO��	x$?��8zR�����t֒�×��P](tqٰ�~VӬZ�V~��-����{���G4�ԋ����,��n~��Bo��N���0'Զ������̑�0���f��
�I������m[y�+�nk��[��|5�#q�;�MhK{��d$�9^����ꔠt>vl��'D�^�.�~�8F�	�[
����$��KQ��K&C�̚L��ɶq?h����ߙ���'#D;��8����{bcP�ڔ�C-��ߪn5Bj��}�W�69l���|�smso|ʡ��y�`�\�m���#��ߥ����F~�^��+Cbؘ�Sa����=��ժ�ZӲU:�p[E�#���ں�>��cģܾ�1�|�VMwE0��ޗ]���zO���0�1� �zu���6�~�NL��E���;M݁���[��-�����=YP	oKރ_�eԙ��{�����m�r�WFN���A(�U �Dhv� v��4��3ըƪ�������`�ԙ�{�������=�� ���������]��o�vtNMz��_�H~�P� (p���[?��{��� �:�!%�����h�)��V	���8�3΁I\�Q�]tC�iyc<�d��-�@����I�����ģ���_����[��"�V��J�Π�b(X���b'��NP%�ayW|/mj�,�tx����VTg5t�48�W�C1�
5,���r��O��B�z�0� �}@�1~������	E��b-�n�'rxT�Z��S�����}aE����8�J�h7�n��T�s�`j�t��N,B�Q�����T�SQ?WR���_�ު�XQ(�r�ZF�_��������έ�L:����1T=?i��M]d�\{IO4���-ڹD;D�v�	���z��u�-}��+�;�=q6�H�0���ߪ��t��!����V�\~-�Pگ7<A��u���
EBlt�'!��/{���}j�2õ,y����42�q;d�q)��� �.8�\<���E�r�	���t~��ZN,�nK��`{xd�Ў�ޭo&��8�L��v��Hy����������?$����n�~2N��V4#a��߾��?l�k�����L��4�n��r��8�&���0 _�N�S��
[�f,����ҺqF�&��D���(��&S�KD16�u0��	/&|�#0@zj���}�s�p��ϙ�FdM�s��Ê�j���6��,�_�g���O���v�*���z��)�y豁����=�-mFx�	{��@V*�	�@����~A8��{N���w9���x�Ճ�<��e �?��^��8;·9g�}�+ò��c�:	qu����}G������/{��1������vҗ�o��k�K_��ip��{�R���ruX������6�eYo��l"t��,��c��#��W �e�&ONم$��!�Φ>۹�.x
��U���;=�?Έ%&!s�>ܲ�x�"���:X,!]�I����@��.[�n\2
����;�`B����+��쿮QD�KZZ�A�A�A�Ρ�n���������;�k��χ�k�f����������@�C���n��G������w�VӵC'ʎT�sf>���}濧���F.[�U����/`�:���?��/�k}Y�����)�D���P�p�#�/�K�v⧿o��OOn"�)L=����F�!z�[x_�1#X���o�y���=��I�Z囦�i�q���+'1����jQv�8�
�!r�ތ�ʠ��)���Ssʮ̕;�d�5�`*�s.�����>!�!�a]yX�8�)g��s�H�w��L������_�B�v��י��-��.�9�����c�]D����?���8sϹف����Y2tAs�xг���`��lgi/ z"��ݸ��W�:E�hۂV�����Np;��Rt��Y��bT-�?��_�`R�/TvT���W΃&jhh0;�6y��>���h%8�BTS��''A���[����ql�kJ�Ā��P���%-�F��"fi��\N��7I?�U�آ-��Zf�.�7�I���Qr�L��#�:6N�y�)�F�eo�C��֓7�������4A��W�ͷS\����w]�_��|�%^��坭1r�2�m�%@Al��I'���h+'bé+R��f�����T�������@M�L�z	Rh����� �x�_n/�,�����R�
��2�vb p�(o���G�b+y����O�w�릟ցu�~�[��/�tE zkuDD��rm=�1k����LV�W�<���x:�hnJZ��Ta��b:�e����WY�
g�UM���`���p(^P-xP�������;g*���rzC�2�;ǳ�3'���Қ������x�:., X+��}�����O��D0*��g]�G6�	�ׯ�^W�fM�aV�IЄ^���m�Z�R
�D^�R{�o���t\26S��95(٨��\ɃP0)���� �eӄ�F�V�{�����o1I�g>j�0�}3
7�1[H�zI�� ͭ$�������J�*�h<���R��;U�"o ���~���=���	u����[��DU�Z�h��)`O��|�@BއK��J�;˟ �}�7}��8�M���N�[o�]�_�@��X���=��Q	�q�%@��Ҧj��,h@���S��]S�x���oR��Z$����(H߂7
�w.¹�Wm��a2�,5*�N��S1�V#���3�jcpvH����k�'�u�
��\Mv��,��y��25��/��ml�F�(�<6�}R (�`,�V���Q;o͝v�^C�v�'���*�jù��y�]*�GZ�`a�����!>�=�7	\�I>�ʿ��C���R۵��R;K���f��9c��F;��?�b���i�h=�w�3҈	�T\)NK��w�Hnb$(�����g�-���<����ȯ� 7i�ę��f�(1Mq�(�Y�ZՔH�o ^��2~�?#�ql���'yLaD�w��5 ���)�Ng�t�n\h��P�s��+�7qf&�_�>k��83ed-�fٱ�b���O�Nɷ��/���z��jۣ���lf�RFi���� =G6_����$����(��)�����A_*���h��B���偆�WX�"�V�/�'fcϞQ<
�,@�������Lj���\~/ioڗ$�����}�`���$.&���԰��B����n��/�M�`*�3��њx!ԃ]�j~�y$����X�T��^�#Iv#��.�ZE���9��
6�0�}Q/k��6��;`���pG��}~i�e���	�v�K�q�lwT���9����{N.Kpħ��?BRI-�z~�[=����/���w?�Ӧ��*K B��������܏��G�xS��Lc����A�eE�X�&9�,yZ��k2n��l=�i���l�� �؋Z�
jx���_6�Eo@��o�HQW(�(k���0�~/j����2+o-yB��`pӎeU�%���͜ho}TE�h��"q\���6�1>�:�K ��S^��Yt���9���� ��6$\շ��D	mg#��a�n�	 �p1 �;g&1�	L^�4+��ť�N׺��c<�f�w��O�9�9���[�D��noX��|٥A����:j��Mh#��U{�	u���.�^���茶� {R@�f	n��,���Q\��fu؍w^(���1�yѱP�s}�l`l��� ��چ��a�I��[�x�,�C|;B�:ȕz��.�jx��[lb�7�3g��l�����C��uH�1�z �)�R��<�Su�{������D6�B?Վ�ϭ��&�����W2�~ ɜ�Ӫ�C�"�=���=�����F�r��ɲ"+Mޫ���5��� 3���Z��Y?�� �̞��7/��c�4�`2��;��ЧZ��$|�hv�ϡ��N����6}'���\��w2�����s2�'�F�q��uTa ���M��V�g/��w-PU 煮�(D�:����è�l}r/̍]o�S���t���1Oԗjgu�� ڜ�u�˷�?�����7I.�Ա�/�������)�߸��Qaٌ^�����B��V�i�h�k�yf$f���6Lk�Ϙ����VG�V�� t��fc��ը�i�������X6Yz��( N�r4.��X��4�.��`���#j&����J�����$: ^���:�7�sZC�ޟ1�w5���H�x��VX�f�����.$O 1�(<�׷���R}]Yr�1���?�*�?����J�.��y��,�{�ư��l��3��qk��(�\Ň�D���^ܰ�����Y_ON�\W�-D��|��1�@��aB��bE�Y��k�}j�]�|��yK��J���x��T�8=�J�%�YS+��r�v�Ȃ3��U�B׫���l]_1w�}"I@9(�#��ߦ��i@���|��1y�[�81��贰kC�v�a7_njk�iWuš���؈'�`9��v�s<n���,֤���r߳����"�����E�V$M@�پuABw�0�e�xcA���!�KM�`5}b�:/���f)�u_~�=��y��3i LV88�w֘Z�X�-�]���.�sq.�=qa�����kI�l�"�4�{���Dv3��UC�WpC�!�z��ҏ�藀�.8�>l�1/��������x�I�2LΠ:��;��a�n�3H��A�@�����ޱ_
��;�,��X�.餜����ܳdO�?Ӕ��	Pd�,����s�������d Y铎��2���C3���A�sW����{J�]Vk����g?�������3Q;���U�0�c;.�ҠΝ9��)@�]Fr���H����-��7��{���w���Pq�����Y����]�~sMI)6U[�QI c��X�V�4:Ē5�;KXxd���� �~$N��-�y����(���h�D�� ���Z>�3�y���m�d���A���$��F�C��������vrE%/i�0�&R��XY�1q������'�v�s�Z=46x$(��������֊�S2n���a��ǲ����dt�h��+l�6X�'�����$z'/$;�H��U�Ȯn��	�QI��(��~�s!�<��]���z�nSX'�u��P��D(좓մ	M�}��
<h�s�M�|�M�-���������C�u��#��c ����B߻4��YS���\��������l��u)��1�m<��i{�SA�1/Z���8�f6g�-�r�͆��gj��ۚ��S������Â?��y6�����B_,��C�u�G���)���8��L~�'��
0,��L0����z���A&	p&����δe��V
lR4f�'�����N��T�qr��{��b�7LiQ_hbK�SV��bi^P�-dP��.۴�7@�z*g�8��9���+�!C[�����Mσ��̫���
�n/���lҨf�>O����ՒܭD�Zp{	Ó�n��Ų9~���5��Qs�h�q���q�m�\)h[�����Z�����Z=���nO!��Z�۾���f��`�D�Ă0%����fy�Vv�h��~R�l��2�����CHE�Eu;��"X��MU�s������ؽ�Ȇmnu&�^����i����ۜ��;qұ���pە�\%��[x���M�XhW��!D�k�7 ]R���h;����g�ߕ	<�R����	ę�1��2G����g��DA��o�����E��^ѕ����E.�vG� �P��}���>�-�J�SoB��>US۱�|�w��U��� ]O������%�ygԨ�y���y�[����$���D�Qt��c,1��B@Oe�+���Ho�[�̎�RXP#����)_�1'���|6��%l*����_^����*1Hц����V��X�n3ިk�{���%	�y�dÁw�0�玳��e����z%������>Ǆֵ
�,e�R�|2�x��?K<܇�N�5�'t����NLG58���ʿX �Rf�����"��B�Ь�����]Ϻ�{N��l��?���̳JP�U�`�9����"VG\��ve)�'͓�c�>]��c�����g>[۵�K~=�u��Y��h94ƒq��k9}�InO:�B��B'�չܷ�;�U��3���܆�s����%��U���el�g���R�0�4g=��:�z������4��4xCx�|9Z'���e�$v ɴ@�@B��6�'���X�f(��\ ��.�N�7rŊ�i_��z�[�=���rMFճ"S�G����n��G�ŕ&4�jT�+�O�U�k(,Ow_��������3(�"A���Z��y��Xe���Υ}��\�����_�N��߯וv 8�;����A� )dA�C��n�D$HR�t�4E]7f��>�x��QU4�oN�}���/�Q�
ߪ�˶-I�M^D��b��Xu-�8jb��Z��i3x�fh����_C��':41Mc'2����KZM0�_�VQ��m�z�%����SK��}���O��ˡ!0T)�"2E)S���p%�z6|w�LZ�T�n�Au���K޶'r�%h�d�ү'o�2�i��=�1�>.��v��aùd�m���f���S����>�����\�i	ʃ �@�a��T�k�.Û�B�^��¿�U�2 1k5֣�h�����z�@}��� F� �I֮���׻�u!L!��aK�Փ����~�![w�kk34�*�kn�9�2G.N�sIG7Ǎ�uM}i\������uU�caK�.$��/�x��ȃ��@��y�;����[��yDyF�K�ܶ<�9G$t�6��ƙ��GI�T�_u^�!�4��W@���w-z�]�H;8�exCa�5)�S17u�>�u!���3���T�B��<�������a,��ޠ��<�Kؿ�u��ۯ�,jͼa��b&3����{4JL�q&aSա�9��쵴>�� T`�w��~�_>��� u>��+^�ј|�hH�{.�S��*ww"p�D��m���;25
���C���[�x17�m$�[��b��i'R	���m��s�X�|�`�ɍA3��@Hhd���4� ^ĵ��No���C��oO��+on����q���x<2c�Cݭ�؛��ug�������Z����ƺ�� B��Jk���J�7̚�M�oFpO	��D��r���.q~[��ą���֕(��Ţ�B��`��F&U���{q�������Rl16�EQ!3�Bį����%�V1�V�L*��V�IpWN�xyHb�Ԧ�o��������p2�t�f�r�hT���f���ԣ�'�U���#U�5�Í)�?���~Z$-�O7x���i�h�\�Z@�-�(m��Y�+�f�uHK�����H������2�X+S��.=�q�E� �"Wb;����v������Go�g|tj^Z!�:=髞���/���g�Ľ�^q��̓�\����I����ξ�2%u\������t_��j������䩻y��\iz��Y�6�c�*�٬�Soj/Iz�Z�
\d_="^�������tP�����"^qizA5�ce�S�������d�+⠖�cÓv1�ejO0����O��`4���8::�����ÆX�l�|��&��zѵ��7K� );԰��_EEV'Dk�����3�X �r���zS''@�;�ŹFT��s�n��Mߣl6_J���B���_K�5�֣�Ԗ���AϿ����V�&oMy�9e<�Դ�֩���qi%Z��ǀ�$	�aU�!C�+F��� �XL!Έހr���B Y��YrC�������l��/�y�ڻ���_D�w�Hl؂���=<�,�^��b�yMm9˗=�䭶�3VSJL��uwB7���CpI��:#e�P��=�|gW����T�"-	K�V�1:7P�q��ܙ���W{�0k�3�60��U	���Δ��F�K�-���'�m�̨g� ���T.N=:�ig}��e�휹Q�-X����z	g�w��0�p��z9���Z��O��m���ƃJ����D�Ky;�>����=44�%z=���-�Y&&�찧�A �k\o��/ѩfGZ�R���/Hya�35�,��E�ڦ�L��+�2G	LoV����l��8��l��5��d����H�l
'�r�e�ZtL�mK@�~pf:�k7#�`�դ��:�M�U5�����&�̗����3�It�`\�E6��sF������f����fx���wws�_��<B�I	�uƌQ]�S�Jڅ/-�4Ui�F�J(�z�����0O$׉�P�_�Tvst���=}N��|d��xml��g�C9��5���!H��܅a�� ۷���y���Z��)$Z��VoTI:��M��1i�d�g��CU=ۓӗ�FR��cJU�������)�coR4{N�9z��R����Yt���h��Y�x۱%]��幜 ~�A�fʇ*�>��c�#zNoSaR۾r�nئ�������������⿲��ir�k�'��P�Еo��O6Z�!��穩r|��1A�5�ep�R{i{!'A� +ER��֝�"�����z7CD��j���k9���7�SR��$�TJ���g|���8��%�x��Ds��-�	^� ��Y��v���i�AH����6X��H�Qr7{l`)9��2/7X�6��L���a�8K�O9�J�(i�	���N��Upe��ŨZl�����������oqՍn��.�f/��78��zSk��\sv����J���gX�Q�Rᖕ�4d�À�M�Ѽ�N:�=&��^,���-���+��>�(y1�w�f���ҥ���G�ή���̙%�-3�yM��P��*đ|���pp�f'�w�.���!������Α��*��d�jހ���_-K�Z�&��p�{ߑ�ʂ��i�>k?١+���`��p}�TT�cq����?�u�n%N�l�w7*�F4M5�b�G�����&��b[!;�B�+���y�I�a���n�H�;i�>3��2��C�� �Kص��k�@�(�6h"P�5�Ya��T}5��3��?H���uN��T���W�ڂ�hu�����)�Ŏ-q�� Y�0,�Ԅgc������y�i�uR��u1�0P�Yy<������.�<���*3��G��=w,��d��n�V3�jZS� mZ�������x�h�^U�W<*��V#��l%=k1P�h���w���9��������o�-y���n�N�ru[������-���X�R����e��R�<�p�Ĺq+�v.{f��J2^�"��A��kC�;�ˮ�^��"�Vn�w���m���������/�ɱ~�8��������h�}�6p�����1+�m<��מv�k�{H��ڭ;`Vo�u (�YQ�R������wk�h���Uy.�s�&�W/w����-��G��~
_�ȹ-U١W���y���ο.�k/�Ϻv>�oS�ۉ�˞�dݛ����B��!�K�P{#6a,��&��a���(z�
?
���j�t�l}�%bl?�R�D}����L�;�׿�;tH����=�~q @�2z��$w[޴ROL���m����@�D�S��7�Ҳ�W�<4�'��C�\b!;�����^��2��L;�pܫ�8bA��`1�k[Ag4���IZ��䣒�ߡH*��^���}	�,CLe���mģ��^�{ǡ��p�l
{K�\X��C��݌ģ���5m�� ו�'�/�f�.dG2LUAu��۱n��xG����!����^IZ��nWB��|Q�L��G{nϕ�>�Og�-�8;�@�<��/����ieU���7��v�/�)0l�\tx����|l���4w��uf7�E�����k��QMK�t�5�ѵe�)���H��R;�0GY�����jo
c�R4�K��$u�jd�f�7%��'�L�u��P���� `�9��l12�r�|*���5�uB5�P��w[Xf��Q)��䊪m��fU��,s]�y˃�т
|�6s�8WV��<B���HXŒ]�m)��A���@�L��������d������\CJ�������A��XBݫ>v��)���.�Հ6rp=C�e!A���c�v��M�^ŦŒ̐C`�2�ߡ0���������ρ��h��sqf�:@#���o�E?9a��Y�>J�ᦍ+��E������ƚ�^R�I3�TO"����,��9XE*J���hk4*:�X�rp_��Z��J��YsQ�>��L�(J�u��B2������^��7b���K]�,Qcٵ?���$GK���K�ԫ��<34%��8�m�'�u~�,��0��s�[��2�J!b.��;_ͩ�d��ie��~����(V��@x;h�����L��.�4]��y̖s^���뾏	+�����0�`�B�|���B��~�?<���NF7�#M�@��%�X�=u�
��#�!��S�J�φp܄_��?A
.5:���ٖ�U�\��cruseM^UF��6�"����$ɬE��Ƕ ��ʁWގ�`��_y�ƞ���KL���-D]�C2:צ�y�*��/���ճ!�F���X�t��t0N��J+<�phLE^�I�-��"���
�>&��ֵ��7����:����=j�j�r��.�nx���Y�	�0�i�_�ٷ��K�-ʕ��ؔKe�Db�V7@\�n��a6gcSO���9�W[���.�<�(�)���p	-CX#�FS*$�d�1L�TJ�c�)_ 1���`��"l�n�&� ߪ�>�Ƚ�rh���M#&V�[b�	��qL��?�Qh�D���*vZ�X�RWd�z&����C�9�f�K�`n�s�nSz�匪J��E����T��Tᤄb��\C
�]7	���%k�%z�O	�NO׀6�6e�N���w�`Y�:J�G����2ra��z\�ynU�z���<Qc�|5!ٮ&/h1*�Kq)�`���?�fy��_pͧ��+�Gq8�~D�.]L�G��dI�m��uZ�bCsg(=����S�R/М��MH�U,�Rf �z8���9������ �$��B��c!��ҞUc�T0�2��\-(���y`�Q�m7X�t3�ig����ƑA���c@MW���)�7ճ+��Sy�$�.��e	qo�{5>	�8e��J@�'��âkn�b�ˋ�J�	_E�5�
��:טp�3��a.X�G/k*�.�B�D�Z�(LA���1'G���]9���I]y9��c�maW�K�3z�Q��/��O��W�����,K4wD-�h�=�L���A�i�	5���g�%&:)���.��)��l�k��D&J˒y�k�+t�ܢiR�_%�p��$V^6A�o.eq���k��
���+Ѱ�Q����r 
���K$,�T �'P_L��|�O���|��,8"�6$�(bT����qk�5��u��0���X/(,IhF�"��
m ��TE���xokU��Z�a�|JPaR#6����G
�	6A^x+ih0����KD(ϥD�X�xvӂN���x@��Lǀ=�@�\�p�n�K[���5ً�\�����X"i�r�:��A���L}���JS�j�����K�{�F��ݘ��]�����_ټ� �1�UTЁ+�����G*-]�����ß�KL�&����!����P<�J������6��P0�e\e-�|�#����I�J,�H�[8̩���A��;[�#�'���3B&�r�ս���o���(.%P�P
 4����׌3�\�ȸ�c�T��B�l(�ҊnX���[��~L��Ю�ZR'&����X�E`���3h�!�ZZ�Qc����ziBGǇ_֯[dj�ˋT:�R��=��YQ�"6�5��4��i�z6&%P*�)�*z,�}1ݫ�fC~� �/غL��pm�1���FT891m�1@��iY�7��a9!܌�J�>քc�$���݃��֜�,U�e��"U��=�φ&� =���T1Q�pQK���ӦD돏�����x~#l�6�����Q�l��d�LOSb�ML+��`�8*ڇx�w��2�o�n�e���ı����+�Cz��v���+�E��w��ΆҴ1�Ig_�����O]�j�n��M	�Њ�1�>�S�ĒOū)��)�Spս%�ԇG�1@�ɼ��"X�r��Z�y�sAx��/X�E6g�
��g�����q���P	$���5�ɗR�\E��1u�Xey׭j�R�`vb^i�ɗ�Ծ��y����s�m\��h:z��6B�(�+p<ؑ��O��]��ku�M'I�/��n�BpY��br�7]�bQ�ɳ�av!s�k������nq�̹%Ϭo!�Qr�qea(����B�ߙ�3�cP8��(�Ƕ%s8��.��t]/{3كXak�s�T�����aҟ���ުVF�ݤQw����c�񪄋}���¹��2>X8����޳�k��� ��	�Ӱ�;�������M�V<z�T�X���_Ɣ��WEM*���E�]�s7�<�E��g�qB�eTW]�=�ی�^z��*&�x���ˮ������6�ޔ۱q��|[���J1��[DgC�{V�(�����~lYv,D%~rGֳ
[x�)�_��l�s�FB8JZ�m�Qפ>p)~��/fF<%��R`�bI����Q�>�Hf�{���꽖��Q�Z���>���6)44��b�UK�dT���4��WtF��5Փ�e��S֮}�����	]QR�iB�X醟��VH�Q-��E~�N��5t[�f��
���ǣ�Z&�'ő��N��8�4���G��w�9��c�e^b\���Tл��.2�M��>4�n���ߩk���	PH��v���c�%�ۨ����i�cn��K��p����%2�����~��@P����C}�bq� Vl4\TO4#��:������KOmئB㳤t;
�<�n���vMg^��C(�r�_�,�����_=�.���BQ�Q˩l6����M��fd�X�5�
,7�N=�2H0���-[�����W^|�7&f�mޔ������irr(�������.��:y\����ܚ'Q��`�/�>����U0}�K^�`d�^���­֒��Hqǟ-Z^,��5��$�w����LR���sG�1��A�Qq�.Ҧy�|
rK�r�B�C_���0��P�7�r^�г�8�ԑ1�{���}��[ŷ������v���M��[(9WBW� k�oύ��o�,l�o�9G�7��&�S�pE#1T�ʒ�q9e�|����,џ2H�)����!��:�G���%���m���B��1����|�3�
��+M���d�if�)��A�e�Hٖ�Hp����*҇����6��hįN7����_�и�4Z��P<�f�E�� �`�OfU���M	�B�^��!p|Yv"��nv���&�5sN��z)�^L��l��B�)3�9j�~�x��q��)|�����̾�Dy�^���o�"�;t���qd��Ѳ��(.��-�Q堰��16�83����M_5k^�_gUsݲʾ��f�8A)�z��q8��2%���=�OK��	o�:�^��-��85q�:}��������l�ӂ\R���Y7�O�+���v ��b�Fиc�g�H9D3l(=���lW���ى�QA�˨��L*i����xĊ�K���LP6O!3N�������cv6���rZ�T�,�������A�\0A*uj3�����f�ce�LA',��8#�A��*��л~ߡ�n2o��W"o,ytY�_9�l{���T�<�Y��e�]����U�k����}��xa�Y��]9L[�]=���O��rɟ�\�<]?��eaM����˹o�@��(���A��^D�z�y�C��%��� %ē6�ٕ�?�Xe�ixk?;�k�xݟ�zLv�w���<=�VL�.l \q���֎e�U#R���@��(���$�L|�٢���Y�ټ�!����	z�
�hOɪ֕�f���Ϝ�0nM���pR�O\�Z��-�RIUj�O�:+�M���9۵)�����54R9���XRR��,?��Є���[kE}���V�-	�P�?�gc�i�4��{���`��p�C#%�\&������]�&o�t)䠻3�F&�g�����������CƧ�[5Z7J*vB����$q�Ϯ&1 �Fiua�	z��f���E@����8q��__b�0\�";t��[��I�M�G*�X����u����L�=42r��s���o�#:�'��M��_!z��c�>��׿'2���7�ᠿ�Y�O;@X���zQ|d�+w�qc�~ˈ�q�f�"�d��vX�Sq����j�d� vy��b,���fdr2���J{��6
��6�x�e��o���M�< ��SŨx�\w�%��~}�(G_�uuj×��������Jl���81?�Q2��Ļ����[M��zhY����jT��U���c�s��~���9�rp�߿$��4X ���ϡ$�
�?yMO`E����dϑ[f��=�Ѳ����6��^�����q{�����Q���QcZ\[�Aކ8��T"�)����\�Wt��N�W�Ĵ4;� ?Dt���"uy��=0�(��׻�pr|����m���4��OW�_L ��RQ �*���a�Z��yض�%c^�q�I�*�N)�����:Z)z�M)��.a�vw}���+ε�h@�N��B$�,�R�7xe%bJc�3�;���p��O��w�<�Ҩ���e2���䠣-�+d�U���U��.�BĢ\���|�N��ĉ9�X !�n����u��+Ue5���s�S}b��j���d�ك.��You�����̈́����<�3eA�����&�r����uT��R%�y��S�l1����؟l��]������V���g��Sꂸ�9g�^�M��	��t^9O�겫����ϧ׀k�y���&�>�Jbf����jں!���A�=��m������'AH��2�
���ƈ}�vT-�����:(g�i������1�ƻ�ѬΣ� $��T�s�~0�X�ƾ[�.��Y�9H�����A�cYH���tn�@U�����K�t.R$�5"���~��J�B��Ø��UY� �ߺ�h�74���͠a��n=�d��	��FOW�-֚��g:Qh����n��`o�G�=�.��H���`�1}�h ���z��7-9&0FTҮ��Љ�;����z��ސnVe&�`fA��a9�T!�-�y���F[�vd�4���,�yd����q�����wĈ�B�*  �=��[��n������k�x[ΚE�RA��d'm]�j�_��^�&1��,$H}O�+�y}]��p�1[+�N������P���αF���T1���ش@�c*��]�S�GteW��6-�o�fTJi�b:�F��+L�ؾ3熀��-��+��t�g�s�O���6�bp�H
r��t���&̕>Z0B�w3��z?}ao�r��Oy��#����^��7��Ǒ<����P�sl5d��n�&�齰��e �7��� �m�F����^Z�\������WHyL��%*Hڻ��"�9�����ϭn?�ߴ��Tx9� g ���E�n��D	�/�c�K;���p��3	9�c�׃�"$�:�R�}̟I��x���^�
zo�3��$��.��9Q�F��h����T\u��M���	�ߣ ���X����IE}~����W
��E�y>uM�^�C#�P��)h;��X�:`�Q��u�P�٪pv��Ǘ���Et����h������`k3�T��B3�J�雨V$�W���H�EI�Hј)h�����q��n
y��:
��<	D�����_x�]
P��t,+Q��:Y�xg(��(��h�q?���F�` -�Z�g`��QC�d��#���)�&��s�������7���ls*
KΘ�6�0�������fR�G��_���ڵ�Z����7���Ǉ�[@A<�y1k��T��;RJ)� �Sz��qAZ�^:����e�C��ٕv_?�'h{hJq��5�V�����W���D�ȓsjμg;֏��äp>eT;�,g�\�w�f��L�n��R@���n�E����J1��JKH�&h&1�\y��;܇S��5n�3�G�q&��F��i�������W@[���A:#"��G{r�X61 R���S�#gNKr������W��	�*�O�{��P-���=H������3,ǩX˟�=���u���,���zm5qX�2�J��;���[ݜEL�o�s�����:���Y�X�ޤRe���Q?�ܮ�5{m0�Q���Я�]�ݙ�-$&s���Bc�3��#�(I��i]3ϝL�gn�����_�����)�m��*��.�6���J���񌹙��U>��i<yOϷ><p�L�����"�����OM�[����d]!��m����6,�'�%�ݙ6�Q�[�D�'?�5Hu�L�!�?mߍ��^�'
׉Qf�ا��������i����|~Ңc�?����PW:	��#:(z�C8��9¶:���j`�Q�J1S�ř0a�/L�at�<x!|�T��9MZ�����1�*3��hy�aYZ��t? [���|G W�>q%e�q:+���ӽ�Մxۇ����x�|~�ha���,1�~O#��/�|J�ұ���蹾���M����1�N�R4��V��]�(�<���}��X����!��<x�[h����c�q	��Kl��F~���=��o�A����5��lB���e���E��5�ɡ�vJX'd��Q\yxs��jqv	[K�:Q�!+)Yw^9#�?g
���?Y��a�%[.$4��S�6�mkU�������Įꆉ�ė�Zb��t��Kֱk310���9�2���uLm�9^�ɖ�4�AkIP&��8��^��X�W�H� 8,B��ʊJ��@	)]�R�����8��(E�\�ة�,sA���➤Gz籝�}�6�u���|��WA}�
�L���b��w��j:�[��?e�ѳ����9}D ���`ɭ���Π�- ���M0�y�2���B��ͼ�x�5�f��폡
}q�����h흽�J2��V��&]�?�\��$:C���g��*����7�����Ą������"o���._�nй�O����O��ap�+5nТ�{ǁrhrUr���K�,���~ԕq5E���dȣ崩%��=����낝8J�Q���!$�=����_�~g�����E����-k@����ٗ��y�^[�01+O�6ᾯ"+en����n�4	�Y�^���	��ں
0q�Gig��[� C�Ϋ*"d�uvb-A�J����J�i�TĂ>��/^Dt"c}��i0�)���Zᘛ�s7?ڇ��mr _&�S�����z���r�*��(��r����؁�dܯA�.Mu~�1��W�1Q���"K��-�yX����.)i^�:���b�=��5� ��y_l�w�U1a��yT-FjBh��{�RbT��id<�x[���b�]9��!���.6ܑ;}%�F�j��VG(�\�������p�Jī̙tF!%��渚&� ��TQ�!1k�����,;Ng&Z�i�2a��|�J%b0?�Mx�y�|�z	3gM:��،�%���E�vaù�B.�[����M([$r
��=���@QG������������/�-���>d�?��su��✥;5�ֽ�A�,�O
S� ]��Wo`�[������;&�eQ���p�Ø���ncŶ���GM��79�*����]��Y�=������,L���|���zA��UB��rc'��?��]���E�P�O_8����Maj�	��N���@N ';ާ�m��,Itwgu��դ�3ף
�����@�'ܫ��Wf`�y`i\[�\1V��	V^���S���*��cB���6�5�����%'���<��Q�Y֪�P����c����[pks�]a�B8w?u�`a��t�(O>��Ê�[�}#�>��.3e[#v$A���tY�j��s� 	la޽G�1�Y�g	���gN�>M`z�;�7
%6��8�\q�V<
޷^r֏�e:���/6Xҳ���6s*L�2��#��<}!�M��ġF��� ��!��Mz�֭zHH�������Z���K�1豾��LW��C�Kd�#eu�����$/�;�qt͏S\)#��\�jJ�&b�*d������!�Ox9��"b��i��I��ܕ�U�=��k=���y/�~ut)^�������n�DLL���2��m���Fp�0M�p�
�i��U ��Jk�h �|]�&a��D1�w���PW��3���?F^܋C��1ՖZ=r޼��b�?�����`�	$�w�]�ww���,�C����݂���;ܵ�s�8����c쇽����YsV��}9|��@�g�X仡�h%L�8��)DPn�D��W�f^�ɳ	 MR�YZ�|����P�'��l���Cz�m3H3��7�19�T� �a��J�#$��5�Bd�����"e*���?w�0*q	?���2,��>���Y�	���P�MS���>Hr���R�n2lA�X7���7��:S��&=��&���?�u�~媍f!؊�l �>���n�'��H�Cv�l�;�!�� ]���7�¥�u��I$C�r��\�t~��{b�/!_�!�jϧ��M��F�4�;q���ʹ���������Oj�w���%_T t�IDi'&Q7 -E��b.�ް�s���#N��X6R@�j&������i��Y҆<�A��X��ٹ=]|hGxa�<v/��3$�!�q��o.b�%
"�2�ʌzR�D��}����G.���W��'����Ѱ����o�����c�!���F&�����������o�fX��;#?A�ߠ�7����kP��	H"���z�Z�1;,}��$i�����p5�a�g=���R"��{5�<�t��s+[�.Ǒ�)<����������9���o9�5g��o:G��V����ZԻGS�͛�,M�/�2���	��ق��Z��S����v�����潿��Y�ߊ�^*Z���������z#�BTouH�ps�� -B��[R0���&y������H�H��q����R�����EՅX�?�Z�j����Q$`�Z��Y��]���Z$âJ�]2d18
C-���Tk*�bX��LL�*)C��Fo��`w�Ucr�2�����]�5��D��2}���6�mxH�B�|�S�[e�#�KS����%W__�D�\���3���'&v�����I�᫲5�� ��Zܳ�t7VD|��%��I9��$d=�n�����s�96O`��嬿�E|J�ݜ?%�O�3�o�k�2���p�(gd|��t���W��0A��훬wKc)*g'y��),f��a��?��CC���FȈ4X~��"�<�,&X|����	5�9����Ha��E	Hl-lX�6�g���⻹sz��ڕ�X�"���=���H?��*d�3��;���ڜ�狒M��3�2v���J%ɲ�?�|�	�������k1�z�#7���qwE�ݠ�G�+� �r���y�ظ��ҋ�\^d�<��"Э�Wk��h��y�x�H��q��"���Bf�5�8�����uF5��[�>���ܟ���ZNP�}Z�C�M �,�0�2#ͱ�J��c�1|�[�o0O����I��o-��\_�j-�wMt���u���uʊlm�WY�Nۺ�#D	O��2Z��8�T���}����!�盥n�o1����>���AS)\���쟊Ԅ�i��l��-]¡��M������0,��2�w���(��
���OI�9@��8�/BZy�k���g�6��AY���Qes�!B���ؕ��~j7Z���F�Z�u�&�E1��n�kJ�\�D(J��	!��i�I����^ܟ�_��{�T��dR���˟���"vj�J�S&��.c�Ŷk�r\d����\nQ�^c��w��IAi#Q� �n�=?U�@�p�o�Y���ƅ!:ؚp�������X�6�v6Hd�#�[����ٔ��0����`��5L��F$�T�d�0�·�h`��M�Zޣ���&_�;w��er�����UZ}���I�s��B�I���2|��OI(�f�M��Sǯ�h}3X��A��j�O�K�N>�Ty�_%�������"0��9�٦�H�����dl���f���@�#o��Wd��{�^��Ɣ�]������;�L�	�M^�Ǩ�D/B��!���)�~���@�?>Wݥ�]��)��+x*��eڋP��>^8��lq���[��&�oS���c�V!�1#�K��8[�E)��t�-;6�'S�EC��RWn������ޙ�Ɖ�#	�kof�u�x�n����=�l͒�^y�B�if�L��wE7_�reՠX'�3���]�7jqX�<��F�c� ������t�{4._�����/k���BDǌW�QQ��+��gm�ōW��������җ�l�yo����~ͺ�^@���T���}:�;���k�h<*Ɗ8B7������~ʫ}qo����Ǣ~���%�z�Ka�;do��T=�!%O�c��#����<����;A��������vU�X��ޭ�xqu�r+> ഭ���lw [ԝ{q>S�?���k+�?Xy�{����7J�	�ń�
T�!]�d�-M���Z1ז���@5�Ւ�9>w+M�� �	w6�f�?��:��^�	��F�6���b���;,����_;����	���N�P��s��E�od!�/ڦ;)����MP��l�9kqK�D��e�t�4;�.�B8�JX�a�~����~\S��5�7�ƥb=@��V��s6۽u��Ü��w��wWO�s���^�	5��%$n�(�A-��bz�h�D� /��g�l�U��'��*���M.)�'"���H��x;/v�Ȑ&�^�v�7�s���I6G��BC5~uf�N��e{�K1^�dܛ�<���13<>Ta�p�	�D
MU��`����0�d�{�,�b������V��y8����?����57���m�`�_�{����ɋ�ԫU
��,��ު5<����A�0�]�I���g8�	�f#��IR��%gyj��������a֝�>��Eޜ�j��Y�6��v�z�|�; N��%B�Af��A�oS��ԇE�s,߆Z U��4� �ݽ3���E�_�T��]�\�?Bbk�:�O�clXR�N�=��*D:�Y�c��t�B�s����tpxx>�_Ͱ����U��/�4whoew���G�6�X }���:AdP.G<���������y�T⏲�a�����Tz3������W-�p��h��´+�}����[�K����n���hj���KO/�5T~YX�^[�٬�Z��	C�ټ�e�}�h���hv�cr/����?
\��� rc���6����+K�����	���P����8F�˚��*A�:ڝ���ǩ+v!4��角q��d�'^��h��˯ƚF��k{&�JK��Ad���,|���p���Ij�۠�z4��Oc�[���9�-�#�.�"�? rIH�es=;�$���IcP��$��bWx{��fٵ�P����g��,櫨�������"-������o�=�Sܝ��*䭕q��(�{��2	�}!z(ZMz����o��V�yu�٤�jD��|�H~�S��ʗ�C:#o�{Y�}9I�P�d˛�� �Ǐ�BP���lY�!GC@!�'��t��e��:�� r��g��}[-��zZa�g�~�d I e���07�Ak�1���$�I�W�EM]���b~�t8۲�"fIB�0�
(�s�un(ם[�s�pZլ���٩�Ƨߧ�}TJ�����c]8�cY�_��h��gc��,���:$nK`��\%cd�3^S?�\xJ��ZCo;��6��K�����q��D#7QW���sP�V�f��|�p��>j���?({��|�AG��؟Z%T�J��8�%e/�:H\j�|ը�Q���5'�9��L}������(��~V�cZ���y9>��o�[V�W�Fw�h�[���Sܵy�?r�3M��&�.H���gN2 �,��w�t����E>�p[�~�P����ŕ}������5`Y���w5}@��\���!�۰���]^�0*T&�3ê� ���g�<u����p�_�Ly�
m$Q��s�
1G8��x����`�z� ��s��/|�^�kI�(�������Ӷ�Zhk߀�f��+����p��F!�+�|�]���
��]"�:�+d8���jE���Z�x��l�Uw���>��E�M�h����>��A5,[� !m4q�i^֓��J�1tYV}���X����L�fpq$[!����@$S�d�P�L��?�5-yy+	E�rB;�"��͐'����>p�w�5r^��F3�i�^&�U�M���?�i����6I�r ��%i�mo�a�^P��Jl�";�s��F-.Ր��ɯa��%�/��X=#��MX����W20K �Y�`���=�b�>צG�t�m���,�5����v疜l��]���I��r%�}ｖ������	� %�V!����x�a�9a( �}u���Y_Eue�X?�r�h�o�x��W�7U�j p�boS�v>�>5�z)qt�YQ�z��:����wXi��h�[z�`��ݝlhB��-���K�����-�G�L�_��wfn3�/�20@L�hq�X5^���}�]h��_���N�@b�P���wCFx n���v�{$G�c�*�f�����*���i j�����Yw�gs�*յ�ӵ1+���D�Ւ�g����q�E6z3���T�!��l��������`��$�$��`�&�o��OK�p���Z���%@�Q���A?�tY�uU�О�u
�����@>�����l���`�Y!�yQ۞˽��KRV�X��������!G�2�N�B��I,z��������vp���>�wh�|@��Iq�ic6q�8�TLZ�8�G]$��슼�'P:�b���ܵE[�Ƚ�x�r|@:���ޖ�C��!+Wj�eHZχ���Ψ)nB�ic>� ��Zimtʝ��		�t�V9I"+<ʿI��(F��%`�4 W�y�iP��Q?�	��62�7��iϽ�������AG�"�R��Y�@�gI�Ԑ~>�=� �빾����*��?C�kk-5p�_��3!G�ΐ|<�#�_�LA%mS޼��������>$isM�V��oWzْ���.�<!��V�B�sʌl�b��S�/Ͳ%[r%�B� v9A����:�B�B�fh<H��T�y偟���bF���NbE�+C4�v�Ϋ���G4��|�2�':0�߿�"��g�Y�ʇF3��ص�T�~/�@wq������$���2��:Ǻ�6�v�H`W��C	P�F�
�xs^��0���� �5�Q-��D�ƚ���}�ǵT��!O��&�y9�������[�pmbQ����#x���I��mbH��P��	���Ω�rd�� mj����μB������-y�F��[J�F�h�u��M�h��N�]���t���'k��a����Ƞ�S�đ]�*�ȑ�.=�w�L��$�<�*�Z8�H�]W+�qX�0�,�l�3�.?�����O����xu���²B�{��"ܭ���JW/h���.اi�QH�ѭW��v���u=8��:��
4�ï�4</=��t����Wm�.��V�7`v�c�Zj���5�x&��4�xM�B�-�����*�����p'5����v�����?�Û�U_��;�vc����Z�ݘP���ϋp��6ߋfux���-�S�	F<唝X����}�h8����Ou�K4,�V^_Z���
	���葱�������y���<�L'����`.g�uz��>Q�o{�ؾ�%���\ys�?�(ʭ�?��Z[yV�We�ma��~@:�ii���
S�|�+���<�4 ������I�m�7�o��Q��N6���S�Z;$7�����H&L)p�\m�i�q�����3�f3�� d6q IY��ǧW��3ش8�`�07�����=�j�ϐ<p32�����}�Kf^t��#�3,|R<�5��F7�a�yp�QHKR��"�"JT�z<�b�Kպ៷Kr���]�m<�Un�}�Z�gis�B��@�)p��)�.��I�>R����'��F��-F��/p&���k5��*%E�C��}�=S�u��e���Ix��"ͼ7�.=�N{.s^�)�t��ng��˩m��	�9�(�?��Y#������D�ޓ j�#�@f�R��;�������
<{uד�y1_w�w��P�j���U��>3��R�)���	��co��m�,��Gm�����Y�i�KW�f��p���$�� t��U�rÿ�MZ��\ң �ɐCX��	��?3���?�B����kPV�b�n�0d�+ �J��6
^6L^2�����Y4'�4�é�x4tY��|,\�~�M�a�2�׈}��|)[�oR�ȟژ�혠�Jtߒ��kWu23�	�Mnj~��֑� ��݅�j�eF�Bא�ocs	0�Z0����� ؏MM�](�� oŮ-S���|Y9���<�������z0�_����V�?���NCag�"L����ʼN"��w���0{tbƫ�b������w�f�?pϛ+
��bãS0e����'�adS��rm�
ŭ=�G �B"7�Q�^mka���B�"��b`&+�)�K��?�Q�W>�^w�2�u�mĳ8RR[⎨��^����!'$�3�>/�[]�F�9��y�=Z�L0C��A���l�a�i���N#�Ɓ�Li�d�⫫�/.S������a/����HO{H���Vq��r�P~��ⷻ;Ĝ���z�k�?Q�McИ̩ȭ�3����-�cH"1W�?[�4*"���Щ�t���۾OM��>�Z�P+Y)�K���Rt�R��X_����q��[zpr;������O�$�OCe�ͳ��+���e���Lv�W�B&��Y
�+\���=�|ǽ~(�<�^�h�A2rxé��;߆��m^�����-�jܜD(�+2��ӠE_s�ũ���{1�m���P�����=ZN��"`�mY��a`��]ǐ��a3�����ov]S�V��1£��w��v��h����j�!a8kr�Wa��`a歨|՜®*��[[�2�|�HAIG�O�N� �D���'���]�YY(P�1 oN��؞*N��mP{�.���Uy����C3��� ��U3_}7"����-J������n�>,��`D񍉻��f|�G9O�<�I��vf��	.�̷� �I[|)W���z��o�w��5�\Sw��9�R��S���D8�D"�'oѵ�a���LR��xi�Z���0H!Q��9˖�����T�;���E9���&�~-��W�]�C 56�]�tn��oz��S% ot���*RԀ�� Q�$9��;w�	!�d�3_��f��}��I�⌀��:+�� {F��d�i�;�� �����_��7U`]X���%ے�9
j	�P(W0�`��z#M�̮}���Q��L�l��7���L�s�=�7�e�G�o�
0|���H�Nv��f�4��~$h�-��n�z��W�Jo֬�Ĥ�X�l:�Sɇ������<O:���*���]o�S�f���g��НT�t�����| �X��5P�
c��,�L�ꅍ�J;�mZVqjE	�3�ē�ܾ�R�`�9�2F'�Ze�]�;!w��ㆷwޕY� ,ɐZ-�|uR�֤���U��
Y�ՄC�,A2V8#o��8��՘]��y�z��d%ǋ�0��W?ڿ�ا����9���D����l5�vA��-��L$��
ϴ��^��/S�\� I#.�# b%����=v����{H.h��c]�Ez�GL��*��3$�h<r�����T�.�>��l(��2���k�Z� Z�����v�p"BZ���,W��p$a��
i�Mv����2~���t��9(w޶��[9�^O[0sm͵>�QW�.p�y^�A�w�����O���7U���h��ߊc+�F�<X��|�=��E�B��S��?S�V�8�@wa�}�X:6g�Y��|S�0$���1�"HҊ"��j�z����Y㬫������{�fL���dF�4��"a�sSV�Κl�ciץ��J�Lyv�պ[g�D��I��Я�p�p ���Qɀp�˄�]�G��4h�Ia1u1�>;��%���n6�
.fW���J��<oMe?�TC�9�5�:	�I��<?��0CJ�2	�E�ZÔÚ��?#.g��]��eu�q�x���g�����筻��&�vͥ��q�mV/���`� �S�ۄ\����|��E��l��haʙ0�����/`N�	�T�?��Z���1��Lg]��,�6��z�"u���5f�
�Q@�z(�I�z�5Un�T��`z����&Wc9���|$8�:s�Ń`��$y�}����0kn������'� m}����l����D-EH��b5,����_�6���eGD� N�T��$�F�=�iS�z�
P����hyr�}�)^3�ʪ�r�c�)Bai����R^�n.ykZ�2�rD�>ѩ�cAu����W�q�7��m*�����M���s߶K�yn�J�GL��=r�g4ZW��r'�� �fnH3\��s&�׆���T����%���Y�~s��(:e�媔@T���qA�Ra�!o��fZ\k@aƤ�f�Gd���r)DF�;�:Ëo�8o9��t�b��=�о�p�ĶQ�R��v�>��N3ҹ���*�좖P�g�
p��O���;ۧ��y�I��W	jӛ�-=\�t�h�l)P]7��w��~��0ԁNP���¾;��{�����j�ƪ�������R*�ӎ�t�o�R���lL�?է���4m���k�뚤-�R~i�7�$��Ӵ����g8h={�N?ܑhܴ��sIH���V��M�V
�+���{JC�sBfst�����(2 ���gj��LՖ��۵�+k>�G�����T�ʗ��5@j�מ�h=г��f��A�K�y`>'���Iǖ�mg":E5qf�j��z�E�0���*�s�V��.p¬���=���Ki`j�,9y��FCan澩��Q#U�J۝_%�<w֯�����P�iz��D�0��^�A��	5�� �2p������ϰ7ڵ���gM�Uz�d��O�ل�R.@�C3�kr�N��"&*:S����8��6q"����Փ�R�`� ��Y-,��v cU�}��K�y��k�E�A��_��XzgN1��K-��]���Ұ�:��<���g�߾X�K�v���B�T,��r�<oPZn8����hb�do���O�sG0^A�_�Z���z��ӞҒgiY�Eߝ�����m����ފaI�/`��c�ƽ�.P|0�K��+btؠ�Nu]�L7�q@E���3�3�ψ�J�;6=�a�д|U�dcǚ�z�&Ua�)�q�<+���̠��mc�pZ
���P:�H���.}�Su�wHk����	ޮ�y/��2<uMGUG��x)[lHm�(��o�e����M��>���D��G�jC�o�Ƶ0*�A��_��2�PI���)kf�3)NG-\��N���v�)���Y��������y�[[;����i�G_}=�,�����*�����ۣ�Au��De����h�Һ��)\��k�CB�]��'):㏳Uo�ı��3K��Z_�8��-I���m��8�y���n5�T	^�D�����J:1ia�j��q�K�ʡ�˹P��F�W!5�ƚ����4�{݂u�`�y��f�OPe	P�+Am�w���a����R�T�vEZ��:2���)��b�Eճ�G:+&ʭ�E '�}g��%e���灁�R+0���Fr�~7]|q-}����s�y�t��r�U&�:�?od��/���.H��'�w>@@��jb{q���f�R��(�-��?[V)A���s
͒�m#$��ri�Qk4�}~�M�ӡ8YｊC�����t��;ȩ�g%�q�ߡ�K�e��N\��A�7c���?�R����Yv�j��z�)����Qj������n+�d�`�2�7<9�O�����+�kx�-_��tŗ4h:�����7�����徣k�\� ����0d7H�*��2��@����;<* �1	�?��:w?���|�\���u�]�z޳�u5�&�/k��A�ɬ0'X'��o�w��v.��PV*��H!��)��K��j>� y$B��'9���XRi�_G��Æ�9��{������t8-5��N7ዏ��C�����)�6y�8�/�$V����tpJ3���_��:�9g�����A��h��?:��R[�O�8]U��톳��$9��^�E����bR1��+g�ݜ���|Y�m�����R���M��ŉ�ʘR�R�7^pR���U�A�tzj����L>��3��T2f�LP}��}�j,�r�~b�|�o�{��&���?��UO�j�ڢ�)��z|�%+-�i�UTSR���3lI�{|��#�X�D��n9B����PYWY�����@L/o�����)-�S�H.��g�yg���W���zl㈌�i���,��%�6��pH n/ܤ�w,{P�I�m|X�uCbּJ��2���.lA��wD��ձ���}_T�-���A���:tt��S4��&m[uV֧�Nu���A�M�"q��g�����l;h2UH�ˇaY��BeU�IƔP�?y�I?�Ń�3[��{�q�S
�����~������4LA��8��z�#��N�+V
�����n:j1.M����%ʀV�*�e��Ƈ��J�k���^>�}�H1Z�S�%��oBX�d���a�{�U8�^3���#�&�A^��؛�N��/�,a�ј8w|0>(�/5bQ|���WKB�U(L�C���ɜB+H� <\FYbݵr����;�U_����[�R�7I�6o�M�����BJ��m�U��'�9�/��X��kb�+�5T�E5��(<�~p��	+�}�Dn"�[���b�N�zc�ΊYv�ڙɛI�,��[���IH�Y�����̢�y�����ޔ��g��*O	�'��z�_뷭$�rJ��)l�	�֔�	&�Zh��js�T���Z<J��أ�D6)�}X7K֣F����מ;��3ũ�-V��4h��o�5slɕ��1�{1�be�"�Ңѷ^t{�t�Z�V�S��X1����Y�m���PY��@]�Ò�yR�q|4�E*���#�MQ�?6�>�F�n�%n����_�n��'] o0��H�8����A ��ؽ�\ˍi4�!>9��ː��BV���G6[$S��Ä3��_�X��n��G�O�Zڗ���B���|!�'C5y�irk@�S)7umУш�u^�>��`YO�A]�"��8�QU�0m�x�}��LTǌ��/�c�-���s����D�81�͗��Y]����gC����Ӡ�D��M�}䓀��S*�Q	��o���̍�Fb|�D�|n����j�a��ϼ�@�^9(_��CQs���OM�o4��Z83�"�E������Gf���lN�,<�C�`���e=G[��L�w�?̕�˅���m2���C���{Վ
��h߮�2=�2�BM��8���cR��lz�� z��f`�ŀ�Ñ��wB����)֡Kq�gL�l��"���U�Ht�������{��:h�|UW������a���=]]TJdg�M�W�j�,\U��ypk�v�}�����M0a�2�'&�� ����%Z�-"IOQc��`� y;���\�>R �-�T��*
��-1��޻��F����T�tx��*Wz��v���t��a~�l7߷U�[���q�O-v&&-.6���X�nY�Sɥ|��R��:���l�N�j?t�ɥ5�'vm4χ���A� /:[�I�9�=��
�/s��O/��DL]c&����KA-i���f�y�bn�{�UR��r�ڙ�%�C>KJ�Y�K�=��z��\�褥�}J�����a�e����ѡv��m-���c �+{��A�ɱ8Q���^S:\z�hz�_g4zё��x�aH���a*�L?���M�c���.y*��7'>N}FP�_C-����Qҹ�W�^�^0�ND�݌>�@���i�F��W�O ��x�$H�f��~���>�G5�H?{ �C�S(%G������٤n�}a���M�����@ӵȯzs����eŭQFFP�~\�;�( X�P!�
d�h_����vd�җrvx��`�	��X���[���GZTK�����UD��.�~��bA��١��Fx��j��@�:�L%��c�����gX�d��MT����I�Mx�!�S�bc��:��x��/&%�z�R��ǜ~���8��.�}0��3�*��Q]Q����롕�i�?(�͞x��p��.�6M�7����i��A���Ov'�[�ࠟ�n���4�56���+�AP=}�c�F�6��כ�"��O`��e1ZKlt_c&��?t�=v��D_mh�FA�Y�U��]�H=7�'�&$���Z*T�w������� �<�H/�IXz�"�15�g͏�%B?�U
��(MܴGaZ�NNP6���+zzY*��[x���nm�<�_G����kt�����*B��o}Rˀ<Q�R�3�m@���$�/���3U����U��p##4������������lMD�$�sX�gS�փ�Ź�]��A�z�+toK7�e&{�����]�~F�d�0��Ι�c\9v�KH+���gU�U��o$�Loa�����4t��1]ϼ(���(�=_��ٺpOHZP0͐���@��A�;H���,��9PR����k��q*D�r3T=��1�k��k�i7?<��ۯ%`� N;�,S%�Ł�Y�ܬ�i�r���bG�A�mCL3���BD�|�<�q`#�W���V>fd懸#���#{J�5�0�s��Kz�Z6�j��s�N"���j�//7�_
���So͓��&��[�b
T"	�^&�"�7IB�Y~���l�\
�O�q=#�����I���O	{�_��I�k�A�ȩ9�b5ĩF$΅���e)s^A���лT���,�h� TdF��*gn�pG�<���;���1[��W�@~Wԝ�^�P�^��D�\ș�%�[���<���փ�̂%\j�J��jk+��q,]'5�#�C%O��a7W�̽���|'��e�y����91�y5��s���~��m���L�RQ F����W���E�����'�S*׳Җ��@��Y6���r�v���?3�V��&���[��JI��P�p����Ђ$׻���]b��қ��F�����y]����l���������T`z����
����#�q�O��<��z��-����t�Ɠ� �
��3j͋)APW�4�'v�ѷ��F�1��mV����EN�)��@���ǟ*�C��h��c�����f�3��[�"�����耠�z�Ԛe�	�>U{9 �@����R�]$��	�xN���rvk%��]�6�U���p<R�^M�Cի�&��O	��S,!nz�T�N��ɴx2eȋ�Z�0�w�����%�)P4�<&���&��=�|R��Z�Lc�9�Ϫ��f��-�p#�/�����< ͱ⚋���0�!��Ixo��H�5�T��K�v���O#������|P��=?���?��o�-Y��4V���LǕ�N"�H�V '?yN��[�������Œ��D6=D_|]o�,�I!�v�`�8���
#��R)��Q���dx��g	��'��c��˷�]x��r���x���A�*�q�OjZK?��c�_�C���H=&\���@�n���}5�H��]_�3|�����-�"�~���*�����[�'�V�b�j�o8�������b,@�6�V(���:����Ei[��հQ`쩥+����Fo��v���jD=��(�$r��S��އ\��⥈�rH���̈́sz���\�1���8@���3+���U�6��B4���� ��t�r�d<����Fw�i���G��#r�/�wN�JXriDH�~�$-���w4�	h8;0�b�c�"$Խ�d�T�=�?!�Y� 2�y�k�� G��%�G��(3	/��UzGvwH��f�s���]��p��G�j g������{��
qi6t�����#qkS^��2q� VQ26P����v����ٴ����~�F���j�7����TLH���Sf��ZDC�1����ag�M���}ǲ�:X��{XAe.I�� �Oz�
0L�G�X)[���6Ǖ��,������G�&��b�*]=�t@w.I�dB!bo]������L�q�mPf
��w(qʼ�?�˪�|P~�)�d�?�Tg�2��j�	+� �	|�з�Q���B�$%�����)�b�Z�����\���R������"�b��;�c�J��	�:L}-F��ܦ�3���21g3�x�2G�6-��Kе�W���zԎ���0����Uszq^.�͛k��8��:��k
��>@��w����Q�q��3���YF�JV���^�r�$�W��9��w�6�pf�����o�E��G�;��R*�9�Id�3�ɛ,�%����A��a6c.�0�ς/��Z�c"?�1p��1���Q1����X��9�J�_xh�h��̏�c�0� �*`s�iE�V�&�5�0M�?0���L �9��t�ݽMn8,-�����=.�/�W���AM�F����Lg��Ct���\2s(D��n�t��|��-�BA$�ٗ��;�1�I���*F�a���uP3ɞՊ�>�R���{�����0��Q<��v\���g�T�֐mK���?p�V�e5��6�і�B�(�i�H�ٗ�V���}qLs���8�,���d��R����	�c�Qj���K��5����h�g��S��"��{v��_gf�P��F�$���~��yw��U�X����:�_SO�݂��Bm��Y�$��˄n�V�m� ���7��}�P��S�sA��gL����K�sˢ�zh�|T�:(#�go"����~*��HN��F��q���!;�V���y�f����(�fIr�Ɵ���vq����.a�4[�y��[���Co�A��HԧIu�}2x�|�$\�oj�O�UZ2*`����
xH}0?"
k�� 1YuK���0K�,f����kz�12`��������[WF|��O�����q�Q���V������^�a~��滞����[��y�/o��-���=���*OM��2��^~�V(�R�07`+-���w������j�N����z�+HB֞zP�����`�m�r���$x~�����Od�au+�khR����n�6��Z�̞����҄(�n�]��%��%������">����^aϊ�u��kL;G�oP�Tj�0lf�E���I��SVS_}T+d3A��j@��̀�l��8���GL�Hi�ƥ���\ƕ�����O��1�����;z`�!
Ƨ�DP8}�*��)��XӴ��fV��m��m|�䫗=w��C��a/4�!�v��gذ~ߎd�j%$X�x��}Cuz���]��Ȃ�/���<2��]����Tz�rfa�L�ޫ�����a;�'<�-"3�n/&tǂ�O��ؿ���ڰ|�lGZ�AH��J&�#�8�_�@�,��t�G �����9]����,$�����C�B�����E�����i�{A��;a������[��%K�+1�����̾����G�t�9zt��v� ��p�+Q�X%b"����gք����%����d�|U��������N�}Aaa�	K����T�V�61'�Η�N�z^U�$�Tb�[�^���:��f;�����Mߺ6s�+���sVx%����R~��j��'�45�Ld�B��w��o�$hyq%^}+��>�-���<X�L�@j7BG�����B�&�W1�ä�`6c���/|����p��0��!0��v^�&�2d؊QOQ>�.��ISտ��`���H�NN*,eO�+L�q3�+��(dW_C�
�|���.:�S�p^w�֔(]��s���̖~}�J{�����;1���SMA&��+;�o���q ���)���)�Jk�B�
��+��v���]�N�34�|q�� �Ȏ���V��:*3�ˇ�I�/�ǹ��H7�O�����|G��赜��P�v8��:k�b����FfW���JR �v"����q��V���ò|��R	k�(󈨤�|�a��8�
mB��vgR��ł����ι+�?��/�ܸs�"��]��,]!-��7uY+�K�.TN^�l� v��	�6(��������p��d��3S�9��1��	O(���҆u�������,@U9�P�X~�=�S=E��K�}1�%g$�{��V9n���n�TE���/�~�P�ג�p�Hf(���Ug(c���u��*�zQ�\�Kt�{zf���r���&�Bx�y9SL&w�y���61{5��v�-I��E����i�hV�)ܶ�~�. <n^������W��c�ܐ��BHW�r��� ����,�;wq�
��,���xם,�:����u��T�[`06M����U�ůEV�)�``�KΉ��XU�ͱ�����p�]+]F���>/:�}i��sLZ���6CJP��!}��k�̥�� f��Z_�Ӭ�M��Z��JʙB��#[&���T7>(d�4��Eyl4.��죦a�R��;w���Q��ZŁΌ�yX��Ņ�S���Sj���`����i�ȶ�>���dz+�ǲ��gv��=ߊvf�=�I�-oM[�G�#�;+�t����U;M_���%�Y8�/}�[;CB�6d��݌?��-��Ŕ��x����5�zI8`,�,1�q�4����L�ؓ'${��V����w�N���x L�ևNw��Gԃ�c�3��U��B�OTOĒҢ~��aIg����e�V�cB��hUEUz/�.yB�ٻh+����0�l6�,��}�޺��T땹���fIY�A�����2�2����͉Έ��6�c�(�-�r4�X����.:��R����a�-����naH�%����-�w����!wi�qk�����~>��xO�z>Q��5/c\�`�p�;V�窌=���-n��i���Z�3�Qn�M�Pܒu�Zo�t|�8��'��M&��}G6J�̐��/�����x��^4��g~�������)�	��v'b���93Ys��.�+ ����	�NϢ�t��x���W+#�cܳU���+�� ��G(,�/�����SM�wr�6	����M+FL_��w��[^ÿ�U�ٚs�>ʸ��
����6��=G2p�uՠ~i��FΈW�b�*�0�\���:GV�*6RI�n9*�v/T�b���b�S�!v���k�87^p�a����`���Hk���	���$l���Zcԣ�į�4|(%�`�&�܁Gڌ�qŜ_�Qt��K?�ߩ惡Bm7�u� �R��3zޒq~Y���Ϝ����L��I��'���^��k��`k�c���k!���>Ҩm��l��U�o�1��iU���O���C�BV���ӝ��T��n8����p��Y�*�Ӛ���ZT�-��y0?��6�\��V�	� ���@��BFu!�/����'
Uv�%����q�K��t��W��]F&���ȉ���n9�]PG��J�U�Ȫ=��޿�3���$@>9���=�!x��pW~��V����oYzoa��`��r���C�Gp4�UR,�8du�.7b⼙��C�������a����&����w@���5n��ҡ��_Q��bF�j�Z]��H\}��aB�U���n�!�I$D		mo�?ӯ7}|R�߃?�	C�/�׳�x�����jU�ցָ����Co<ێ��oړ���J`kߔ�0���-�VG�b5�+T�5���K��r�{t�;�S}wU�hJ������-w�O��r�,�u��6��[�������o�z���D�2��vdQ锅�G4����Ʋmb�_�S'�9����@�@y�`�i���$~׏[{G�lKJB��E��D���EK��6P|�^�r�v߯�f��c�q3M��Q��!�U)!����Z��H��GA��G(�.�&CO{nd��-]��~��eK"�����)@9ߢ�b��F`�Æ����سS��;��*S鈓B|��Wce�!��/�|�\�,��kz�w�B�:k|0Mt@��AℏEu��K	 �8^���E��.��| ��KՆ�չ(ћs�˓#��v�\N���w�u�<�l�_ψ���cj�bV�#���Va��]-��Y����F��ّ��\ww�D��x����8�=���M?v�@����T����OV�� �������$Q<r�[:�JU�\4q�[��e�68�~���4!����M��|E��F/��-�=-���X"k�ϒs��ޭ��+��?v"�\��8�����s%��<#��`RZ�Kΐ� [J�Z�U��`�����L=]�ss�?�fpo�����㣌�Z��bp4Eh��BڜEp�4R�LG����{~�0J���m/��_��X�cğ\P��M>#[m�iE�O�}���K>W�w\8���J�g���!���}����Q��q)�����E�5�E͢�µ��u5W��CD���/ױ�zjt]ӈ�8�bF?���׸sX$ e���.)�)kF���MV���H�d���dI��'A�^�P�9q�z�'��topp�mM1�yg�p7��.���U�Ǥ���9t�.F�	U���5Ⱦ`A �	�a6wk��50��vw���V��(��Z�!���&㿦�W�]`y��q`x�iγ���zz�\^�(���S���[�5�T��dC�ײ$i�|���nk�߳�%ϧ ��;˝�ErY*��Ü�-��
\`�f�x���l$٩>�@-u��`�V��E֑�F=�)8��W�V����c�����@�!6�����A!�fk�p�2�����or���6G��L�����\%f�k���/�>� n&y�+���,�&Q���պig���`�t� �͚�t��zE�ᑖiN�>Ć�M� �]�6�C,R7�9ݣ��l�>ޫݒ!��Ea�W�0�v�*�Ҋ@�6����$�:K�&�� 5��� ���DB�Vk�;
��	V�+�p��	5�R[��A���7�z	� xˎm.�e�L�a<�% B�Z>���~��̔t�(��MC����X���q��^�gm1Dr>=LCϪ����-��i"�f�S�9sC��\4+�ӻ[����P�SQ����7�Ï�R�di����&�KY���[��\���ٓ]q����}��J*��qI��.��0�F^��u���pmΦ��������>O�qwn��qq�1��U?�1�P[�+��a,�.	�v�Ċe�?�~����P��"�+��u�S�v��㭙,C2՜��|1y�C��l�{zµ�?X�.dǤ��hX��)��B�8UɌH���=B$֋�-זږ��7��b�d�y5���ҵ�� {�줙}�'8��ֽ|�'�_�6��C��\����h��N�z���8~�?��C�/�����L���0W�hxI����Q�3�3}C㍛���&��RM֓ڛoM4�eL��*�p��lx޸sgk�D�lZ�oR˗���C��M{|*�
�v4��@N\��fQ4G��p��߁֛>$�|o=�������(}�$�Q���2�����}np]yյHT�i�ٷ^���qF~�I+�"�Bgy �/�mL�{��!�uO��7&�=���� 8]u?��`�<f>m`�����?��E�R2�wz'��_b27�z߿nq�<��=�;�T�3mQ?��A�LYF�^���:?
(�Mo��L�4�bC���`�Q�i�	8����g0�8�d%�{<�ĘM�#�v�a�<n�{ ^g�������� T׫(<-�dG�+I�Rh"T���-�)B%C�1���֦!�d���D[�������_���,��Y��􀵕0�ыࡱ�Э~�s�_��B����y&�VΔ ���X,��f�����gX�ｪ�[ga��4�م5�HO�-i�E1��j����[���D�����c/���h��t�*ľd�d���z��+�;;�ą��m{3�p	��:8�i��wv�V䓿��K�O��s�H	⍨bP��g'������4��y�"����&V�$�e_�����H��T����և4y�f�n�ۢ� ����3ɘ��j.��o�� ����xK+�
+f����L4O�|�T����y��Ɉ���>�x%���͌A��6���!$E�ѥ�$��ލ=���L�КځۖS���;	1i`��88�KW�ߖawS��j��=^&��NA�i��q~/�����ˋ�{-+�ƛ/X ��D�U�e��!������k���0�5�?�L4ۮ�H�:�'d�՗ds���uݹ��)7'د��C��k���Ց��*�i����\2��zd��P�1MzT�#yޣ�p�i�r�J'�A��Z�]SD��1t�Ł�?t%�������Q n�X�Y��Z߶_�[��\5�ԥ6��<3ɨ�.a�V�+@A����7F[!boL!�ٶB��� ����
:����SuI�v���>�o���Dt?3�7�~���'��t�FŐ��ˉ��fiJ?uɣ0���'�UG-��y�r*y����}��se�����M�ȳ��݄9 ����/_tW ou]� ��fI��,?uI�����Wb���i�`e�l�`(��u=��UO�g�V�4C���k3��N�hl���<#�N�h�i9��=��vH&r�ɒ�17`I�	�,"o#����C���30?��1��G+��+���rm�"�Y�_�Xa�)�yӚ�U��G�Ӊ!?v�c���6*�Q����`�� '���F���0^˩!<�����A�*!��^_��X�� D����r��w#�ݔ�n`4��]�<���(���f�{��[��%ZS�cɝw�ڣ�����|����*_�m�\���o&�i�yc�ٹq��k=��)*�g4�jeɷ�N�6���
�nm��c�z�St�p��w	:��G���q���h�����s�����Ju��F�i'W`��Mխl����:�R�ܬ����ʸI�%����%������8H�S�+T�lߤ���Z3�=7E�1��?����B�ӄ �0�y�ۇ6lj��3���������Nfx��T�%K�>��2Z��1E�_"	(����]����&[�'�R&8є��k���Ó��?Լt�N��p�:&��!�\%n�<�&�`�K����:�F�6P+c�\�oLt;OD���#qNg����RK*�˦�6�@3��3�n���g�}�U�[M���	�PÈWè�'�K�G����<��sUՁ�
�����#���$�i�9Ə;,D���eS�)}_���A�_��Us9��6�+A�Z����-�٥~��G�0�}��ȍ�(��GK�`?|� ������zT��zXXۀ
���|���inL<�V��+6~K+i,�G���i��Χ�r�"
Dc�H���b��G�d@R�?"󉰸1q,�},�1��P�}�&S�҇>ex;q� `G�c��=�[֩�	1�7�Em��e�1y�o+�n'�l�q�4.�fH�c�$�l���FRa�h:I��Ns�:HN��xpj���~�0"�����[��^䱅����Ԯ|lʞ��T�`= ��l�%=:�R�e�l���
���SaÉ����5��k
AP���v�%Ng�7%Hȶ�˓o��|�N�O�� �
�mD�*X��-ӽ�pO���Y__T��9���B/;Z�WU��g&��4�v�Y�ׁǜK��c�-�+�aU��ʍ�n���=�p�����eh�T���7I+,t�n�������ʤ���9YSt�5���x�8o�(�k�����1��o)J��쓊��čܗ<p�Ss��b�
��A9��K&x��-I��\Cw��ZZR>X?�Hjݤ�ծ;�y�a$�#���� ��Ni��Չ�U����x�g)�>�V��Wވ=�AfT[������Y}�?C���3ݧ�%Yo��Ĭ���I��I�1g"�ʑw���3"���>����;yS�����1�*��J�$�1܎�]���U>)����N�Uu�����\.D�#����,b6�6�-8���,2�ho[��������M]6eҋA͔����u+P>y+T3�?k<.��1H�|����%�R����1�*�%#�ʹ�,	�Ǚn"fK��2E60y�\�>k~/���C�e��!�\~�����\}���i+yE9�|9>
(x�����!�߱s-�1�;W��wƸ�z+�8��Ĵ]wZ �G��9C�=6S^�<5S��U�>�@�HO.��V�X��<JD ���|י��}D�ަ�RxϏ������8A|�������'���S�A9��q�2/($%y��VF�]�E��:�d���`Z��4SYɿ9+�>�'ɞ��nƫ�1ll���>q�.�}G�Q��ߥl)����k���̼����n����$��)�xR����P
��VX��G���jE^�ߟ���z����u�T���aYݧ�.��풫1U�����)�(��s��f���������J�������F��m*����õB����XC��kn�����t�ՇG�t��	�)��c���y��0�ZjG�R�oō�����(Sz��=�=�m?'(A󶲈`?���sYjsa.�r�U ���&}��S�otɢ�M��H5u�l���ٯ5�!ř�B�3�r��ɴ[��֘0�Ϳ����P�a��z�=�\�X\V<�;�ẛ�'��Kw	�����r_�X!�"\|�M��	~�ۢ�.��p����5ԃ9���z|��^k)j��u: ���f�R*�;PV� �!�u(���Y�r�_C@O�x����e�5�(X��I�M�E,�N���P�)k"�0�"�ҷŉJ6,�¹��/3��g��s�x������BKqN?��q��!6�q���:��Z��um��!�U%$��F�o� M^�_Ӈ��y��Y�:�c��j��,�p�^*9��V��P
�ʃ�1"�s�- 4B�u�Y�L��ѕƿ_yY�Ve���;A)��
���Q���3�/��#Y��S����G��$�6����&��*49��������Ts%:�K�����r�*�/A*>����.��@)W�.���݇�i���A?���W�Gє�YI�?q6��]�]��hC�ݞ<���f9��$�qH����q��ϊr�4պ����`h�6���{������^��|h����1 ����;��K������<O��c�q��J��k%�Zg���q�!E������/v�b�	AA��p�ȳ�x8v��b�����v0 ���z���V��~��%W����B��,��{~���%l�sC�.1ι�
5��t��" �P�Fxs��`R��&	�gO����Թ<ثΈ$϶i����o�MYl�Ę�i�o��2�zב�c9՗��x�=���Ϟ�Sռ�8��xӾ�Rێ�T�����Vg0n�?�q��~6]��w+��W���\�_u��Ң��?��|��M��~����c�O���㞭ZW�����r�64�N+,�ZaK�r�8������U"���yPG�Y{���U�FE��g��ީUR�w�B'����i0�s8v�/51*T)�`��g����}�����I��y�y�,_٩��3Yaw=W�f�4>6W��~-8�lb1���� (*���CP��k\j��H@��.[�	2�N�(L��_�K��i�C��I�5�����س�jP�6��$���iU3^������"�\�z<F�W�ZT���H+:�'W�p-��H�)Q����Q�����+ BQ��~!k94����� �������=];t%ϞV�]��d��~.K���UmkAq�^K�b$��9�〇|@�����:��
&�q�������k��`%���_�8�֎����QW���2a�2���^��|��~T�j/�P4��/iJ&(:����)Ҵ���o�j>S�q�4^�_��a�x՞�~�'�I��ޏ�T47��L[*8J1%4�@��b i�Q���R� g^4+��9R�5��<%X��ZgT����ΙY�C��
@��_Y�<��x�}�M	,w`�-ʗ���P���gO�bn�{��&F�Y)*g#���c�ٗ����#�{�����>����ב�T�}�������`���"5-k����ǆ	����(�A����&�+B/�<�
(�X�}��Jv6��X\��;�H�������!����������/5�"�n7E_L�� ��;{�_��uo/�E���a�o����(z��������a����M��iKy�S���3���s���c����-e��~���Saʩ�D�g<� �>�u(���%�UO �b���� ږ�@h�w�Y����n���g\.��2<��L6�	�Kx���j_��ރ^���F_���<����c�$c�Mfr����`�g��g���P�ݔ�����D )��B���HV��Fp=m@NS5�d)�M��k�ˬ�%w ;!1|O1x�����Dj�������v�<n ����WI�4�$A%W�$Jof�u�=@�J^�i�^�t�E= �� �������ʇh�.�3$��0K�,Y�
�h���1񘑊�dj�j�D3�n˟ٱ8Qފ�0�ʕ*��p���{��h���3�]4�B�q�wK��M����K������Ƿ�,�~��Z�ǻ Ux�Ro�0'��|¦%R;{�n�=K��I �㗲�aoQ�|@'�#_F���X��[���#aǪõ~>#,%��o�p����-��f�F'}�N_K��X�\E_�7��Bk�t`٘�G�]~9ۙi��.�!F!\@�p�c:I��M�ɩ��;8���H��	��,�r�:�S��Ko��)���'"|@�^Q�A�G���	?��\���X�ȭ�,*�P�)<�}����z5����x�h�=�!���W[N�/n�b_<�= ���)���K�P�&#d�@�WSf�J^t��M{��a3e�>�������S��-O�C�["�`�x��4p�����
Q�
�U��1t�9��g���Z;L}1H��J�oE����l�.��k���]؋7k'��H/�� ��9��5���:��p���;_f����k���W��&,��c��_=k Q�=�$b3:���Xi����o��r��$�v{zs�`G�Vb��E�_�4�7���W���M��ws�^'z��<`�NX�L8��+;ȕ�J5�/gp49ɽ=n�zʺ1jI�,ę�|�� Ð<��.�q���_;+h�H?'QV��WƓeyN��:��G��\k���	%��1Kv2yʔ��Ů/1%H�u��h)�D?��S�f�N]�&!,���{(� 	�>d���nS�^�Σz������Cn:7����\sqꯍ�.�v5�ة�&�Ӡg��d5��}�����b&y��-�=��Y��{���_u`۝���­9��!o�?�P�(5�1	�/��
��Yݏ�Jq�$�WU�N��U�A���X�@�"x�'Be�V͜"������b �2�`��f`Q�6�g�o��sn��*���	xv� �,�Y�[�we��/f���E#�h2q��p�P̟�k�h1W�=[�ڡ�����'���#I�$����s����R�͍�8�XuƷ��3����F���n@-�=��1�?��jp�;&·���q��ư�;{v���5z<�;�K����Z�F��A4�8+��q�)v������^
�zT�h�8�b��y��EKs����i9�6���sQa� �|���>�~���e�ғ���L��ԯ�Ü:X��U,p��|h�(6��n-���,���v^�Yh�@�w��-�}�������|���h����=n��<�X; �����Q�m��1� }Om��{�7���&~�	�)3Z���=�]�o+��W*�?����u� Z������ue�fw���F�u���k�oؑ�4q�mUl��{����Ա�"��ER#Z��M��P'YZ?,��:�bʞVDB��#Js��	�TR�ܦ��-]	(����k��N{U����^�6��0��O#�����X���&8靰ADt���=�cF5$��v�;����-���|;n���xd�����
�2������Ϝ1�����TJ��L�u�����*�e��
�w��f��01���5��I�w���;�u2W�M�F����(&�n���9U�! �[S��h��Xj�=���0fv(�q�v�ԣ�n�m5���Qno�*&��R 0V�A����l��\�/Z��$����B��ⷀ�P���*(.DE��X0�Rr�Ɋ�X��W,hsF��t�麼f#��(C}Es4JЃ�T��ç$Z�t)��(O����Mic��䇮顒�����Q��Z-��	�����P��װ	��9�K����t)��Y�ރ�V��wg��P�ag�h�4���ɻă�Z�R|�?v���Se�C�����$�b�)�9V���?�����i�����g/P'�>��o/-�Y�+�m�ۚ��hD��4�8�>���
�ݥ�h�YB F�	�gәV�T�oq,:N
��b��1�%�ǉ7���e�CK���
������Fla�L�}:����!4_Qĺ��7uQ���ƣ4K CPO�iu�c�$n'@�"��+M���U��'xX4��I-��(�d�ϒ*�����9]"}�XȻ�`3s���
�ã�:Q���B�QY�ǧ�q��|t�xW�4u֢�ŬT��l�R�ޤ7�E=��-��V��.em���"��y�!4���;p+��Ɍ_g����>(Jؑ�پ�_�K簛4_?)�rU ��W�0�[+�o��rJ��`H����f��2�'����+Q�X6z;�F$ �Xf���aa35n��������
�"Y|���肴~V�I��!v��(@=L�l��D�s�Ŋ�ˣD�2VΆwvW�G� �/OJ�agÃb�t;�(?�]� �v�۩�5�؈3B�;@��/�>�� *G)	J%�^^�.��6Q��m� 7:����>m��̛Kq��3 >��󨿩�YV�֣S	^�v�RU�w��9����x7e��b��h�>R���.���C�ӳ�e�3Y��=����V�K�&�6�7/$�\���j���	W8���ͨ*����M����/yQ:KNv�r�W.��&�l����Rzą�=yTN�LV�qܠ��d뛜H5ߴ|'�b�/��Kq�Ʉ�Dya���N�W���ef�{{4Dz��\��[:!�"2��~���N�̖0�/8���Y�hHB���7O�17r�:k�t�� �n@��k�E
�Y�S�/-5:�@8����Ԡ�Vo~�y�C�Jщ���v}i���!�hy{=��"����LW��fx͡�L-���Q�i�GhtV�	��t����ă
�����G���X�Y�O� �Rb�����bk�l��,&b�� �c�`K�˂�qO����a#�ʖ~��W�;/��~�d��牨�O2*���C��$��q���n�_9p<��u���3.�����p@gB_.�h�HI�p�>�Y�W/x��1ky=�-IH���w�E�MA�?f9h�x���0��㥜�gM���O�~��?�'�H����NT��0��ғp���MJ G�â=~N���!�D������b����96OX�=����Ś���G �Z2�9�q���˘=R�}l��!4|[��
[�vX)OZ�}2�J�M-+>���_1�1�ɵ��X$�ڗE�M��p��a"Ȭ��v�զ�z�=&�p;�4��׍r8�\<pƔb��7|O|D�5����5�ҬF�Gq�X���<��2WS��+��x^�ɾs7��@�rv�#�QӘ�X<�x���W�TN��d4�P��I^R���Y.)�/|
��de���Ȯ�f'���ўE�;$��e^�
��w	Ư�8P��)wy��Pi

HU��1��I�`n���Tڼ�⌃���B����e�6'>���7���T*#���+^������Rj��Pb!l��!���d�\a!���g���2��&��Q�b9��v1���Q�[�i�ݳ��x�O&=6[9K�{,6�#��|�d"_�[�}V�,@Vj�Yǥ����^�H�Σ�-r�Z9��ή�p�8v} �^��}�un�ڄ�;��4���D�����z B={�����R�y4�=������/M�@��^�{��th�;�xm���6H��) ��:�}�
��PS����1F�<߲�X74���{R��ṯ 3���r.�Mu�> će��C>Ӗ28����L��zP�à[i_�Z3����9���y��xV�IwA�EB�����o�m��Bt3��U��t";/�/=ưt�N���8�h��v�&�>�A,p�#�mQj�a����i��5M�P�!1|����x3��,3�|�_x�����*E�2F�g��n=��_���fw�\�D�L���7���ӿ�Q��`C7�a�?*\���Yxr0w�H�9 qT��_&q�cūb#�J�i� �j��k�Q@���6BH��3a����h��v���Ѕ���,CL���QMb�ڡ��GaѤ�|����u�G�@�fmmpE~ϥ�ۻo3׀\m�m��©3��w���� �ɟ>*��Qa��������s���<�%OpC^��?�\��r�
��s@��t��%�ݕ��&��4���dʥ�٭	�|�Ѧ��_�'}�&�z?�br�UX>vu�A��k�ԃ�=Zb��K����y�O�n��������t�. �\_�/�5Ɂ�A�s��2f��@�k]�����y	��Pƭ{��"t;��%h�hV`�56����Cr��� 1��G�E֓泮&.e>�0��dX˔:�ԣǂ�`��������zW��L�,��d�k��V~&�U����j�b0kR��=�?�k4t	��d"Rq�;���å��]�i/����K�[��H]�1d?�����YyXm�t�rs��@�FO��t�U�����h+j�Rn{����Mh�I�F��<���<!h#G�-v����8E諤�U}�{5|E��!���)�^?���-b�,I��:��@1�8a�D�wz��&����:-�o��|�H>W3�.�!�6?Ŧ{���w���������ܧ�S��M:�v��@�?O���ûx$9�X���j��A���K���M?�"��o5��ﲿ���p>��bЏ-�g��'��wAȳ�:�Cē�(�&�?���2�GG��?q�i���#}�ҍz��<\��m�1u�+o�ubO^c;�� �Px���C�TZ?[�m�2��"�<0-R��n�3h��ݹ& �ő٢Kb�ܫ���7Ք�M��>�7�>�d,���cj눔�Swٿ㸇"
0>��̎�xۋ+�~5V߳��@4�g}V82&�i'~���xg�Qj��j�aT�A@C��oh���]8��FC)�x7$"],)?V��	�3�i��z�ҾW~WQ��w����/�݉�r����վ����Yө:CwI��Oz���z�W/���)� Ǥ�`M�b���9�+��^��w���-�V�͆FMgÚ�U3�������t��E)��̺(0*d9��8�_{��i7c
ղ9I1�v�@���d��w�	����{�t|�g���!�=���3���tC\���h��!LHQ?tS7�$�~������4�ua]�_�Ȩ�L;��i��9��/C�7'��O"�$f����.F���~^�x�z�~�Th�:1��J��w2�X�ɷ�,?�q~[�����-�\~�R'�[��a�b���}e�2���LKp\�X1�"�.��ַY7�b�v*�Q���zg8�p�"�����B���H���k=�:o~������l���|�1��t��Ʒ��ދq�z�SV<��w,��M\⤗+�\��75t�j4ƻf$�g�N!�վ��A�'�6���p�ó��g�#4�����˧]/��<-��}ag��VFNB������e�Q5M�o��o^f�(@�᛼��w�Dx���y�m�ӱ�Y,�mΞ��M�O��bc�M35�}�S�؟��>�߃��-�˞-�Z�������%��:���ݼF�b2Kp�L�����$�L��z����S2u5�k'��U��yo�"Np�*"�N
+�+ ���J���'�aU�n�f@�1|>�X���������7��t�g��ZVo?��Mh�r�r�;8��<Y �I����v�m[����媴&..e;���N���w�
��!S��c��LC���lzSL��e��q\�}��IԨY��X��N����&2�mk���o�6��
��������i�7���}\�U�Z�]�
�Y�C�>��t����M����%�	[D�6���@�0жdS��iu~g���x�����5��3>)���^7���a���rt&T���Đ���X���2��o���N$�����NS1]�P�f���TH�5����=���R�5��˓��L!H?���f�`��x��Uܘ��0����5�= �=�V���C�*���(� %��/?87�}ypR�j��v���!�:��>�݄;B��E�@�Wn��f!*r/�sۦ�҄\���aκG���g�^��m4eqp|�^?�h�7���8
�O�괜 Uu��,\J�e�o҉4ǩF�s�q�>��l3+û,\֛3�w�	�c���{��n��8�L��O�2�R����z�0ƳSOH�'��%�l����j$�ǲ�r� �Ӷ��ҋ�B����?�AݾB�Ѩsg����7�m;�v�Ĥ��L���c��������fK�yr���}:Y{����@��w�[[�,�Zr�W�>2�B�3�������i�̬,k�{�!V�j��g19 ��ׂ�+��jm�L2�Ӥ��F8a�/9/��dO����i�,bե>�W��a�fw޵��I�fQD�ޜg�19�kSP|$��բE��Yc��4�vJaXw�J��}��"�R��XPP Rօ:=]��
���n}��_W��Ŕl�:��c%h9.W[��z��o�$�:A�s-]�ˌ����2��"'�v?y#��:ᒧS@�1�/��U�ǵq'��iw�M�*���muמ'�ZN��Os�q�l�ڊ��eD�B�[7��Z_U�J�#��R:�ҫ�K���U���3g��dw�!��hq9u�'R�S��{<3l��
���?�M��:��n9�X���撅�Xm�kjL����������҆�$s��{�p�$�����	8�è��F��C���{��8t4�3�ኗS�	�v:�.��!|>W�ՎG�2v�v����OW��dt��|ĉ�2�?�ZM�!������h��h��E")�����T�RZ��Dǉ�yd�#N}�NjA+��<ͷ�3!E��D�t/G����u�\��j��!�B�|09p�N�RԢMn� s;��v������F0���.9X�A�k�>�ӚO�T1U��z0I�cY��J�����ڴW�
�L�s�/7^�#����gK*<�&l��Y;�V����j�5�l#nq���s4��Ǭ8Xl��l.�li	_Mm�eY���n�b���=)�������N���6f�{8nV>����L3$\�?ɢě���YM4���`9�+�x�?%�p���F�tO�#�TU��Ʒ[ˇ���ӟ�&�\[m�� .k$���}[��#��1�l��tfח�Л^��<����.%*�>./��}g-����`҂�Y�-^:���jBiv�顬a󹩡���w��Y�5�\�S�J]j���z�,��1�c�t�SO�L�5ŕ���{/GY�Ry�۳Y�$�)݁�9��Y�fuLbM���Λ���z޺y�pv�L���ѫ>�����%�Y.?��6��ˉ`P��n�I8�6l���>_��˩�p^}�����D)ת�%5��9��!"���Z	,\k՟_c�a��Gsr��m��4��.�L��:򁄪J2��```��v)PtH�S�ʬ;��,?Y<�e�4��LBb�ן���/�s�v�TOtY�	U^����9���eB�ȝ�E{7j�nX�����--����2�{m����e��t\� �A�㹨N�9<K��&��ګ'0�Z�ס�.GY�d`6�*�^ewG��꽷��E�i	��NWܙ}���)��
cA:�
�X-�H/'cd�V;��Q��^�q(WϺ���a]�����@	f<�J�
]�/�MOA�SҦ���>��v?��s�@e(v��������7y�L2*X���k����a��;�n]��b���U$�F���̟~`��|���\jU���?� ��]E���Z�V�M<6����"��h3�iqd��t�"�C��]��*���\x$���	����%���Ͻ��RgL/9@��RK�}Ɵ���]��<�eБN/,�y?.o?v�^����!��Xri����'���,������P.'od���~>2���3��^����Sf���)ǆh.⾝�F:%+��Ye#z�2�sKw��f�8�5�ʷ�C���0X��Y��ʰ	�b��Wb̢	AR����*��y\��!��/eh%�:���v��/%锉hְ$�k+g
C?cεK���7��ϫ�f�ݴ�"�˰00Q�ʐ�sbnQ?�S�D��a1��5� 6B��ӝ��3pi5�u�5f���������f���M��$��@4
(��-%�$���L
��Zj��	�9[��A[��?d�׏^�<�P���E=?A����G!��r�+�,"�865���g�ۢ4�O ��^i@��G�$%Vzyh�OШ���b��l,�RV�1>���,��e@8���s�}�LV��\�S�1�niw���1�����������}#�щkȳ=m��0���9,��8WR�(�s�D+���}���`�+��ȑ��W�����R��z���J�K�Է���H����A�ź��A�Q�*��O:��;�bs�����'��'$�Z�U�%Kų�u�H�ʼ���8�@
�����#�xSjY*y���Kܫ�2	��~.ACR�llޣb��맃w�gO���V�������KC񉪄kD$>��N���N> *�>U����r�%�q�]b���ݣNMM
'#�3��״��u�ژ��R�6��"j '�;��ۃ�ʹ,���m�N͌숶T���o�1*�$C׾���՝�2>ʪt%�|d^z�9C�ya/}4�#WqQ�\�57Oi�U�jP���������W:�J������O��q"�R* �(p:�-�$(��!��ĦIX�'|����g� 9����)�Rjb�s\i):�?� "g?�:�漜��.g�k�����hFw��z6�f1���g���b�nq��zJwXC,�uw*���*��.+�C��3ήǧ�vݲ�x�Hr��q���MrpWY��d���=7�wk�Zxhg?���Z�T�����JH����f�u��_'��8�-���^G8���������a�~+t�>�åP��6C�׾��zp�._9͛����]�7�Hͼ�'��S^P�H�h��#��I�Ƨ�"�M!Y�	�9�s��i;�#&�םҲ~����A~����D�����#��F�o�Av�i���`xP�����^QMuQ(�bJ��T�KU�NB�H�A���4齓��"�k �*-�H	����������g��s��e����gm-����e��{>�w*�U ^��Y,^��}�٧PN�϶<�swg#���d�-��6^�3}���֢��d�j�L"��t��e�uv#:�D��8���x55�#�d�����c_|-��ǘ����q�M���Br��,k,���w��<���m�t�E��^(�_���;*	';�Mll#�m�^E�k��#j��c��DC�Y^C���[J�'�k���O�$�F�u�<�䢣�p��+�4�%ǒ��3�����y���/X�C !|������5������3v��A�	~�gv�q�S�Z#�msט�Y!A�g� ֶ�Y�F$ޭ-�`��T�Z[�۳��8�ޝX#�+wP���"g�BI�-vO���n��m�?b�z9�I�G����bt�ϵ�C�R�"1H̘q���P|{g���1��<�B�Zf
"��#��.f.2�#qh��#�ك�����������o����
�O��ƣ��^�>�����}|x�+��5��%�)JMe��
��{��Euqh��i�ʽ��[B<C}�߄Qi�V���Ҵ���o}��}R)������nŦ��9V����K#��Xe�������\��3��}��,������C37�x�<�1� ��w�Y����$g?A�CeƁ�FB]ܺ�%�~N5�k�#��Շ�/���'��$:ϡW���n\��2�&].�r�<�o� ��ɏs��^���J	/^xL���f���Gk� �3O��߀�E�:�_����{W4�:�"3R�"��5O���C4�����7l���p��2����@��nQӯ\MSc�9�/�d��]%����8��ۢ�j`p�`�E-�ˮ���؀}ld�9�?Ʒ|���;��T[�*r��2�����~$ղ߁�^3s{P�!��n���ZF=V��P�5�q�M{E/��WK���
��I��E��ī?�E`7N�����B����c�^����!u��{���㑰�3�K�#�|��ۓ!�9v��n��<����13r�k�< ��aT?�T�}M��j���T�l�C�^+��E�J�?{�ԃ2�d)/�cmt����:�}���λ���Nz��(�"f+p�v�Ǭ��4h�}�&6R!�1��ۊ}@Uw�s��f���JI�FKcE�6.F�Xۺ�^<��lu��J��;��e�������+u�Z����Pa�
��	�P���>HRTn�(�(sVL[�4����a��Y�l��q� ���:�o��L�t~9�!.K~qD�d�������0� �a��F����{���X�+�/e���(S&�٣r/ڠ]pHd��lw��>#�<Z�_��.�K�h��P�����?�y���`�H��)���/a�H\y8�����l%�,�sW���I�O���[-{z���6�EA� .ܝT�a��wh uN|���v��P�z%��x����1�)@'����<s��\�}}� q��G�20�4��*�Q��X�ME_\�=3�����Sb�>���C6e����4����ќ1�{�/������f��y��F�7�;+��ٹ(���u�|�_�H��vܳО3��Cr6z��=����+u��x>�Ȑ��T�~�'�Өs����DpV4�= ���x��}A���Ρ6��D�qrw����X�t^�o.�h�טm)�X�8���,(�AW�a�q#�Cs�b��Z	E�7���AJRx �g�'�=��<����bE�rKZ'7Lۺ�|�\5��4���6�����%��bPR9�������@�D� ��ȉr����/lrf�8����唖��Ґ�aT��r�%�ұ I��C>>��L��̀ZmN��T���w/�������r�vKS�E!�>m��W@���q�͞������>Sk1�4�A�3�d��ڜ{J����ogD*���X�������S�wj�.h�[��������ۇax��A���f%�I�
�ۛ��	b��ݟ�M�I�Q�w��_r�c��C��/8���3b������~��9�H�)� �^m�̀�K���\"�2�;+LQo�]x�Z?+�@���E n R?w>U\k׉��Z��\�a��ff�Ka��9&&{X]W� �N^����!����4ݘ�%�>�Jb�T͹M(B��]H�3�ɛ|��I϶�BM����O|�$*�g���6�C�� ��gƈ���Y�Q�Pp���]�xD*<%� ��R6�;�s-��UEθ�\Q�B�o�O��8j�<3ݓGXv�g��P߽`,Pt�����NscϬz���<��K�W���C�CI���U��o�v�A-�񛨏}P�X�@v[�̳��^|a-�G�ZKl����M?l�%��$=n.�	��w�D�Nem�`��j�@�7x��>�W�c�Z�X���2.II�IE�Ǟ�U�_r�C��]Vra�&&��'�d��ڕ�E���S�cle��0�M�ҙ:�zq���� �[&>�����;��ej0�(K���k�վ��ۗ�sM�9~�6��ڰ�%fF���fI}y�˴��`��%E����������g��� %�/{<�d��6��S���w,V�'�ɵ�p�Þ�{��@`�f�?��<2y������ct���Ns�ư�t5d'L
l��a$x�Ɣ�*���'\��^�tAb����o�:Ck�X�{2:@,1��_�*pӷ�����"�؇����'�==��0�\ڊW��<
ۭk,�\��	�B���z���6=c\��l��ֈYh�T�[馠��K �j�������V�)ێ"���Ot<����qt�ԙ�,TO/�7ς����Y������oo�!ȟu[u�� \p�4������3b�>F�k�Ac�g��������=�%���<���M����W ��.-tmT��^m?�>���5@=�3���j���z����>����C&��	��:?��=�`����c�����%jp�;6����VI7}E�ϖ�΁H�H��Z�Y��� PU��9�̚r�+���'�3<��N�]v\�G���� �5ۥ�i@v���w�w�� N�� BϬ���<�x�e�Dv�@�>MN�kV>�/�D(h�s��~>���Vi���Z?�x�֢)%���*���|4Gn"SE*�AjzG����ڻ�Y���W5�_u<��>����r�훍�8��u~N����;��8^*�6w(*h�g�t�4@�,%�0k��$����73ոb��Y�Ow09�_�
�@`7��#��%㎯j��h��B�ir��;E�)���$���=�:Vn,�0�?ŷy.�L�?��_L8i��T������%33L�YO::�)�k�^�������k3�N�)���8��^0��^Ӈmc���M�W;�q��摈]+j�g��}��=�{�wKi@��E�L�J��-��6��鯌�X����	A]�������_vpp��k�9�.Om1��|opA�9d&MvPS�u�"̋=S���~��i�<ֹ�vRe���e�}(����0��O虜f�%�&�"ߺ��ĕdm��h������u>�y�K��ۄ��G?I��I��������|�cRf�5r�+�R��L=b	-eEӓ\���^�)?"�ӫgx�Ămr:��v㳔0���b�-o�_�
�������=��w/�C�I��q =�*�L�ʳ�|<2���\?�r2���k���^�	���[�s�Lf��% 'v~�joь�²��H?z�[���7.L�$`
\�����f1���O�W�5�����"��h�麑m�~��3�~��\�f�<���HQ��Й��Lw��V�$�}7$cPD����v�u���&Pn�M�h��Ybh{�ۄh����3$�7�+ж��������mI�����D��_�8h�8��ք�V$�ط��%���0�qY{'��F�U��	2�.��:kƑq"`�]g��i�
�N�ϬڊJ@��5 ۓ�F^WW0�l͔\����Q�Ԇd�����㘺����� �b:/�`%���mns0]��Jz2��ӹ�bgP^Y��9I�\+�]�NG�pL!��Y.��b�t����ڻ�:�]j"䀱O�>h\h<�
P�b���̅�g�������=s[����?:u�2�
���S��X�15D���F�0*���Wf��:ě�>yy]��>581{���%}�>G7���c~�;�������_ �����E�e�̄~�]��yto����x���u�#D�6;ۼ��Pܾ��]�
��~Lλ�Ѳ�1�5tN5�Ǘ"��`�S�*-��\����;i�2���;�R��B�lI�`�z��+���	�s��!{�F�h�9D�(��D5>�Vz�CO�<�${��ā�ւ�a�o�^�$�ߘ����Fs_5�[��`����TP�7,��{���q��$�y��6Z���\���=h#�J� �\�2$uy�&26��Up>�7�+��b@x��}8v��DP�[�tm�����p�3�	b��>�� �t�Y�31�)�a�6�G�{ �<8a5\1��R�D�ѣ�+��}�ힿ��)��p��򮘺T��	ʰ���^rb �ІW�b���>��%o`�`�E������%}�1��A�ԩA�J�Z��	����^�XV�����)@.0r)$��#�aoS9d��� ����l0%�R��B�^�m��(e->>B��A�}[�)#�:@Z�S�1m��Ux[�?s��������{<����I�9~oV9im�l��r�����j�]�Hh^������O��(s6g<^o��[�xҀ^F���Т�fƙ���Af��r�ǃ�~;��
dNu�y�rb�bu���U�T�����Y�}a�>�8���ʓ3Ir��(����Q��8��y�T�� ��t��p�٭����@�j��iS���h��ڒ�l �Y���O0���AJ/���o*���b\�=��S<Ӹ��nd������c�Csq� �'�u���/��f{u9��)�c�}�0�/6�����\�������0Spl�2�4>y'���(0�]��b,�g����I�1��'������u�Eϧ߄��<a����1$¯�2����4�Q7|�_c��.��1Y��/w��ԣng����f�L�\��C�~pcJz}2���_���BL�.%5��5 `Ď�ٖ춱�4r�M>e�����
UZ�� ����'<�����%^
h�����5��`�Zg�:�sP<����zu�p�[Uv ��7�ݫ��� ��p<���S��	��jq"yj��a<G���J� X��۸dd��S�rh�׊W�������#��^��x2�}��B��>�姮J�9����O��R5yH8ly!i47ߴU��(���c�?��]i�S�q����n��?�R^�'��0��{�Ɲ5EH�D��=	/ķ����vCv�� � p��H+�A����kxct��/k��(����|��#��>�[&W����(��`~���gA��BL��|k}�u*J�l�ڋ)ټ'��e�dkD<Bbh�	U�BuZb-��-�ZWG�Y�/�$8�������Ё����1��~y|4��q[�4
��sS�{%p���\*׌ˠ�չ#�a�$���Ȗ\�K����І��ų�A��ꛯ��F|��t����J�-͠��=�Lx#�\�D�w��[����m�a�o}�����W�]��\�mɣf�~y�μ��X}g�"����,�|�`�*�0�[-�a��A���d_��X�;�+V�u�:nbx�� �2�['��d����_F�U�o�EK��#N��>��5Hw��qJdB��:�R3Z*�0�k����푤O��Gڌ��d"c��g��@4��of�>ϊ�28�f�*�:5��S� �F^��Eq���p$Sq�m�4���Y�i�G2,�f�`m��[Ͷ����{�$�v&�GJ�����n�i
c�]���(�|rJ���^e��mL����>���A2�Mr8)�+��iD&G�)J^r�d}�}�C	�t���}F�fB�c��7<��3^�E��k�C;�?�!zSO�"�Avނ�<q�9�Pi����g�@xg��J��R�ӆc�����Z���j?���#̪鸑
9��,��W"�G�2۾��&��b���%��:1&81ئ��q�f&Y��dS��1�Ƭ�!عR�@��|�1������=9��l7��rK I���/K�Y�1԰��r9��a�%R��尥j1��`��8���m,��X���u	M�_����i)�O�x��r�HO~I?������\��da����3=-�=���v��W A�I���N��8�8�����ETjʵ�{��Ɩ��g9m�lx4�8 �ݻZ���w��qߐn�M\�hJt���ޘu�hs��=Z&;?�������`��}�vA5҆}&WTp�Ǭ\θF��������Q+��c���'����x�W�o9]j}��x�����	A1�xx¾fy��yַ�U^��,�܅K�����h׎�z>6&I~(���)�"a��c ʳ�t���10�fn�%.��(��|/�JY��}լ�w9��a$α5A��i��I'����n�8H�<�^�\mc#��Ss�7Z6�E���-�i�P�/m�\h�膟�i���hTʫI/�q�*Q�H;�14�7!8M1_TٸR@DмXϜ��7������æ�e�j���ݙ�/� �Oa��'�:��-g�l�vv����ɀ�ܨ鮱�$2ǃq��	���(�p��\��s;9�4gͽ�:�/6�V��?��+��X�l�@1���e��Yj��iv���:K(,�|ab/7�6Њ������'z�|3��~}�CP���h��k��F��_�����)��>��Ĵ��=`���n�䍾U�
=g��>�%/{r�#����
�a�N�)���n��c]r���HHǥ��0�Ә'���/�#�mߤ��G������`/�F}��1�������}���쩗��ئ�ט��C�i�BΔnP��9o��8-S@�}��4Z3��;�s�K��{T�Rrޑ{�aj񁉥#��Py���I�d�0��d�mo�H-+�%�np�U��,P+��Ԋ��^B�+�/$|��������0��w!8C3�s�79CM/!�nOՒ_���m�����;i�����9_��ˑ��� �6��r�*J�0�ZRa�����TT��?�� o�S��Bz�	=%�n^9�V��Cgڶٜc"��L/C�`���0���"���7~��^�Eu�~e���x�.a�;�~���>�� �mG�]Ǜ;����;%��0���B��X%mw���6�Mfǩ,���L�T��ZiT�G�MbL�Nӯ	)�0�8!����.Zb��?��]�h�!��>��mSXm��1&� [��x��n��, ͥ�&�*y��]�s�P����/sK"����K;�?���af�v9V�Q���=�a�$fnX��d��k}��[��q�c'�9���sV��=̻:[b�\&���ݝZD��&{F���v_�v����-NSɧ=ZzOѣ �_��|66��n�ޟ���l��8
��M w�A����prF����
�a�>�f�Ɩ���Z�;2'��%M��-�x"Y�ݒ����& H�Ew�`��"��Ha>dߏΔ�=p�/T���~��>u��^����[T#"��$@��je�V�7��s�vĊ4����g!��:�4v���`�^����7�| ��6D�Y.���M1��ı�7&��3�ű�kA c�Ƚ>_e�o�eϳ�9+�$�3��3R��,Z����s��/��ǰ9������=�Ƅ��x��]ܼ8���l�ނǅ_�ޏ��xz˶�]
Φ�悯u&�y�@��Cݺ~~�E�x�c�Y��\-�4�_S���b�,�m<����ʳ2�.����h
KL:.�:?%y!7��`}}��T�1�&X��z(�H!vCр��y���=Q� ]j��ܭ&��j:&0�9ss6ޱU��
�;��j�w�(�W�|kBR�<+�^���1{6�&��}�V_ZS�*�pW�/$��]	�ң�Ic���E�C��&Sm�!/(���Fc��Wi&w�̬y i�0N�Bł��.YǓ�jܼ���$B|�G��c�����������B�l�q���v}��� �}�0jM���h����a��~�n�Zs���ŲR����a���z���7%�嚼������ǯm�Sv:������Ę$�Ѩ��ׂ�Ӎ���@�}s1ʷ'gW%ͦ E�o�!4ۏ�(�chyq�c~�����ńS��~��!���kLWa�ʦ�7<h�0�Bk���T&|婒�4�c6��wAE����p���Z�����hOCbM-�w,�����Y��M��'c�T�R�ȵ��V:+��}���NƳ�I'b�0��o�ĳC|�E~�1��g�dJ�P�-��{�UHj���g�b��l�1~�Q�Z�N�ѣJ�f���ĳK�??t�&�	F�����������>�f���-�E�J�xk_5�����*���ۙ�y���Gc��dꓼ��~�+/)X�E���E��zІ�k����!��ZgWML��@�{?;Q����P'�'8R�y%��S�t��Nϗ�2+�c6ڒ��-Wa ��V���W���VR	�@��_FB^�I�)�W���A���T��!��\�rquE�GiCT���r@�O��V�ƺl������Br*��1[�*q�=	���tN�c��)y˩W�,',�}�����J&�����������o��
�M)��P%��䈣#*f�}Fn꧎5��15j�����lwFHb��'m�a�RA��cI�\�Ã��Q�/ܮ���c�u�9ב�ݾ"��͕[�����&�S<B���m�k�zy:�B�GE/1�u.�4��K��I�
B���K6�q���.t�ƛ{Tjf��e���Xج�<qz��pײq@�[p��~	 49T�XԑLa�x;O��h�r�D�9���hO+�7Iv��րjL ~�ë4��ƥϋ[��ǵ�
W��y92gm�b
��W �髢A�u�Q��8c��5�
��@)����/e�F��ۛAw�A;o�`9����]
0�џ��5G��v(-�������ʆ�%��+-eŊ���6<�#_2���D7W��*��_(�~�nGX���&;+3�I���S������*/�^M��/KAn_�����"��v�9��>i�G��0�
eg>VpL�����O�v|�"̒-w )�����\�਺�J}�t�Y���՛������N=A����2�8�z0?oꤎL`8�kjR���R����A��6B��Nӷ$o?�m����N3��=�ӂdu_o��$�W#V���f������J##�4����V�9}��9^ZA�{���ɟ���%S�T�˭��Ll��vN��b p��L����d�-��0� ��Co��������ZK�ѳ9�����4�Ҍ[�};��[��?~=�aO��k��8e�k�y �A�[fY@�VCxH��^��O�%�� ����̲�"�z*�XK���wи�1049Y�`@�|��ބ<	僌��E�" ��'g���&�n�*���v�G �ϗ��C)�W��ĔL��g�냫m���%T$��8`�{�ῧ?�5������Vֿ����<��r�A�̖�T
�Ә���W����s�%x�������B86�Ti�H��9���u�|�X�/ɸ�/85<���ri�8�%a����ٗ7�m����p�I6A_���r��>s��	3�'�>�m������� ��I���W���!���~c��^��nE-fȜ�����}��NEJ�xf�^��ޒ%<\����џ����L-�S7_z�3�Ȥ*�;^~�������>�ż6�k�F�Z��\��(F&
�������'�5�Dj ܲulN��	Iky&9J|�k���S
OH"����A�IZټD[g�x���C����_��Qq`�p^�\�����j�6	"~B��C����SvުԕA�H��X�AbF�<�����A2�����u>w�Kݛ�Q���}C�e�����,�}𡉙�ǴNS����R�
��`�lj�W��s�yx���s����qJ��zx�]AC�D����fԭ ��4�(ȉ~+����zn&�
$C��0�� _xT��A�ז3�9�n��Fk��U�&����<�z$x�T8����T��8�oZ��}��-��Ȯ{�E%K{j��G0>��+������Dԩ�BYO(�ئTϣs1�38Ȳ=���\x���5��ў�W�	�o7�P�#1��X�0Y�C��uG��|� o�<�_%����ܕ���A��뮟��o��7�[�9����>���6��҈����'3�>��/u@�U,:����$�"?�Ժ`-��s�Ee�$��g�8�i��?�m3u����a@�����|i��`�*�����7��� �]����x8���;	E��Y��*�M�Y

<�d7	��@ni04��ǀ�|�����r�{|��rwU����v��wӴ�s�ev�̖������L��8�"�2�l-�����E#?��D��e�ԍ��=�6��N��W
}�Tq����Ώl�g��=Z1L���x�����R=�"@eeͪ�d����u^ud�2�Pp>D�,�A�0\%��E����(;�F-�����l�L�hg�6x��T��m7ә{��4������Ɋl�}����)��7��2��&ӳۧ���|�=�B4����%�h������ӫ+��zf	ˋq�}n�P;��=}m��8�s���	�
S�2MA������`3�$�Zq���;�y����F�ۊ�"V��ۍ?~,QZa>�vZHn���{�$kǼ�GV���@vW"�h'�����K�#�g��i9h��!��`A�bE�Zج��M	{�o;L�����-�sإ���*oq��/'i�}��*�����up����I*K[.C��Y��=r~��+�R F��q5�/�� �S���	>{��Ζ �K��ܽˎ�5,5.o��"})�v,�@�c��D�;.qA�A�vɟۥ灟iTv���q��,���V�l>��/������_|/^�
����#tI��	�lV�B�g���s�6/�F�]_�w�Is@vx\��6�g�*���++o�vl9>���\�F�9�HM�;��Ѓ %��O�<=�{.\B� �.`d0����|�H����H�8���6��[(Ռpv8�$U����,���҄�G���%�뽑�s�����\�<1{}D{P�R~>�zb�[&��߶�@��l73(��� ��Rw�'����~����"X���_W	V3�zaF8@}8�kkrxP�k�t^ً8ي�fA?Ǎ������Q�;����0��D�>6�b�ad�>M�k����L��)Sʻ���1��P��_�+�؛��쑸���D���{^Vd��Yʼm�½�v��*�R�q[�,�%��.��92��i��脺��ک�q)<�<T j�}��ۤM�O���������r�q7����Jg���8H�g���"���YZ��z�<ߍ��}�T���0���%+e�T��nc�/`��#��MɃ7GO�$k�=f\��Mh�ӧi2/��:��7�)i�9;�g�1��ںQ�'�A�̓�j�m�Q�3AzF����Z��l�B��g���٣�E�Բ�7�F�U�~���Yo��H���{g_�/G۳oYT���uz3�J$y���l��X�GQ�y�4�)±9s��`���N�����ۣ���~+�\��U���0�����%���ԧ��A�i���!!��L�Yi�)~���gB�L��������JފbEM�7�Eǯ�Y��|�\c���1�ӝ��\g�
K��>��y
� U��$Xae�Ol(`���"��퀈q�z���m�T"5/4�<���_ҚLٸ-�m��;�J ���&VL|�!}3h�������V��U3[3��,WЯ����sk�1h��J ��D&��=�E[!��^:�u.�ɛ�\@�|C�%Я�Պ�+��qbv��J�v�Φ���zɂE�Yʊ�Y�o�t�f�|�h|T^Vg��w.f�p��K[���p�kw��u*
e&lr�F��KDa�p�|hn�\�1M}љ�����P�;�����Յ������M�����Y[���̂�i��7ˡ問�h}g��}�f�`�&����1�T�91�84�=�|<mgd��ٕ�����}E�yw���kI�	�XB��+�u����	g��؋ 6N�~D�6&��p�BC��\�����5s���$�
���O��H��R��䌪�K�i��~��4C�.*�a�5�"�@����#�����@��h�8��Rw54!$e��w�%<��s�4=��"@p��Ǥ�D�Ahra�p:G��]$�a~3)��K���N��
�δ���4��d�i��Y�ք�݂^(����nK�]���ӇXRM�}h������Tf%�E=<*a�����N�X�~�7����7�uY��s�{lo%��ߍ�����y�;ڣ1}}D��Z���e��t��1`^h���KE(�_�On��������FQI����
=������	�Iın�\�����/�|p������9mQ	�ն�
I	��u��T���O��D�k�zW�S���6�$.���C6J�������}�A�t��㦣�3�R�yN���Rv�\��'������Z�gJ��`�
�ْ�G0�����NP�nO}����-j�w�a�<5bȸ	:AGg�����m4mƽ:(��E���t�. R }�lL��`�濅~I� 76�$��:�W4����X{��;r��8���&k���v�y=_�[ٮ��`n>���'��5t�>�3��h�"#�y1���-(-�k;���B!�/U=0�26���X����o����3��G�)k�s��zl�P�x׭�z�=�7�����&��/
��(�b����dĪ�ʄ�Gu�.�����
�q�^*뚚n�+�����w�	�4���K鵽��#|�F�x�՚���A�K�ѡ�&g���j#�:����VW���U����r�F�b��k�N��Y���t�D�r"$��J�OTȪr f��%?�bB)o�"/��`��$сp���+�6�˷9��L���D�)S�iݷ��Hk@�
�E�TO��y���'�}
��n�R�$�KW.~�y�
�:���3R��:&�� �;/:�@}���8.��P^R�|��1VqN]�>����g�=�v�d�����1��TL�=rYm<]���XS�F`��l�V7���^i��I���	�Nܻۡ���wen�xn����,�/�693�<�h����&r�s&��Y2���-��ivl�ƞ5���[����C���������X݂�${M���F#,��e�u���vz��e��/+�N���&�ŀ4�Y@��P|tr�v�V��\�����P��q�	2*�^	Wm�i2�^ë�:OQ5�E��ݳ�:V�V�kI��G"��)�`?����� �6�����ꭋs�H:�[ޅ�F8�\ A!��}]����I�c�Q�#.��t��h�Z�������@���{q<�=�?�]���/�^v�i+|t�3u��*>F�V����N��?��3)ţk������������k��K�[
K��(���-�@|e����g�q��I�s�К�㡍lV���'�t�K�d��2��JJ���?�5�GU-g�^�D�n$ɭ�m���;����+���{��w
�k ��n�����$����h��]6		��'1�n�t��#��1[>h����pdA�=�Y9�H��\�M��f��$�G"�g$a��>�(�!'�f�P�f�|O'L���<fC����e��,
�k9<	��чڛƸ�A��{.����8dW�)?Q(���~>}$f�����ϐcmr����VxJ~� 	ݰ�H��_�қ�|R%yq鿡�_�t�2pi�z�C+�}kP(�U��A����z��r'�9��-a(4>����0^��eϷe�����QbL�H�5EϠ���ǖ|�6����=~~�	|/�fC��kE)0ߵ}9v��h7٦�]��۝fZ� s}��n�}�reZJ����ZЫ�-n)+E=���#f ��	(���_�Ta;����5���3rҕ#}+�/`�A�se��,݋���\�愃�э�����h��&�7"Rh|�}����Cx�z7GK>�#	�<�B�5�������VnIG��o\��^]^�N�Hp�Gu1�˂D��|~}]�cI��g�$��b�E�*ɯ��:%���Q�C�NP��D�g�0WϣK�����!%��koK� 5��Xa~�N���E�m���x����Xӿ����$o��A���wT}M��jAt��Dm�G���p����0Ug���T������`l��ۦ��q5|.&�3�,��S?e�Ҝ1Y3�������xL\�
˹���7u5^1,J%�ڎ�,ڭR��n��|MpQ3U�}M��e�K߈�%��A�:e5���\��V�s^�W�I��X�<d�O��#eo�,⫓q~s�� �˞3Q%����/L� ��'t� '�I�@�x��_y$���%�rg&�U�|ɸ�<�I�w+frD��3Q��D���&g���ǜY6�j�ߟN����.��w�6?�\���e�4��7�˹�<r��h����2���ʗ�����~�Cbp�&�rp��S�Ӫ�t�<��|�(T*ԝ���CR�rRޭfw�M
?4ѝH��M$&��0��9�ҨuPp�אK3o؍�D������J�k�]�pkz�u��Jq:�L[��\f^O�OE��&a���j��%����C�g��B���XUa��:�}3b�|k�Ŏ6ݡ�5�k���)Q��|�["v@��� (�2��	��K������wl�Mc�B�+�?6[�鏿�~J��g`H�.}��ǧ��b4�	ɹ�z�Dw`=�����֬a�,(�8P�8;��Y�:Ÿ<�,�4%.�r�Zc@��{;js�B�����3-e�F�ˎ���[�
/ (�螰N�Q�vv�����|�MI:��QE�V���Q)M��/�2ZI����r����Е5����m�8��I::�q��bb&�o= 0X��?�n��x@�r��qSL�<vi����ݐM���?rǪe>��{���hCG']tyZn�TQe���y|���urD��G#�Nt�j����~��A������I�}U��m*���,t4��T�������5K$�`1��^�������d?�K6�ǿ����#6�Ӱ-�CN�4���p��%$�CT�B���_L���{�14�H@�>�x����_�܎�Gk�;�P��Mp�8O������r|P���nc��S2�)m���?ױ���jS^7Iz�M�Y4{lI��v��ڈϫF)w"�qe[��߇t�_��&UH����k{�aC����D ZйLz��˩L\��@9����_����F�'��x��«�\�q���tt����o�2;��xawvge��h��R��m�5n��/q<RI�i�ߵ9��KKx��S��~�����?q���~X��e~8;����-7�y��1��?����~c�raه{1`ɓ��N����i��AG/'؍���3���]|��.�S��*���!���hT����켛z��_K�i_��o�2�ss�t���T> f������Q�ng���m_����n�s�3�=t������������~ +��l_�f��wV��(�#���N�<�&S���;:�Lw����y���P�
$��`.X��S����[�W�ׅ�˜��_J@-&�p|���~����=T��Ѫ����wD�ʭ��oD��<��_&��X,]���;=�������.>�~F�|���n����k'��<.���u��7	&V�:����Q\���5�6'v�U>�G� �SG'��m��+3)�	�搓����<|D�~TtF���GB�nk0}�,[�a�)��l�������t7.�_����L֘ �ԇ���a�"E���d�3s(�7 �`���K[�sjsy�d�h�w�|������5~t���4;Hz��X���y��1��H^����ƚvB���L��ݵ�3��{�.#|�z�so~W����"/�<u�7��wyd3L�ƞ6�#��M� ��� ��U��b8=���s�o��{'�����/ ��C'G�t������&~����cv�3��Կ�Q4�(��q��� ����}Sv�;-�t=� @�w�k��A�Ѩ����!/l�$#��;��O}��;Uб,��մ5F���5�%��,���N֗�	(�?�~�F=!�>j��{��h�[+����'ϕG{���ty�s�M0{��=��0J�ȬYGo����Y@h����5!�&�.�=�h+��x����r뵥	�$I�M�ʤP:��5�#y'o0��~~~�"Ndj��ȯ���*�(���|B�qNa����'�	�:*8�p���րA���g���R�D�d��ۻn��Z�9$�-���M,���HB�2OFB2_H�Y]�����\�zݍ6��uJ���A��K2��>�Rr^]�6."�@�TB�u���/4~�$·�a�!�;~T�@7��0X�m̷>�n> ��7p,U���A���,�9���umw�eMAA`��oi*���x�]��:�D'�pk^����pJ@��������'exj�ܰ��Z`D�WܒOe�9�������-�_.k���/xYH�ǫ5�W���W�y����1b���/�����I����C�[�5����C�Mp�(""%���%%�1b�(�Ғ����1)�́�h��=?�߃��������]q��+�����t���O�ڵ
�I������"N�u ���g)~لT�p����t�?�������H���~�{n�V�%�v�/�Ѣ�o�R��=����`5�s-�Z�X�=C|o�2�������0�X�<Y|�(Z���#�z��_K�듳Y�0��k��vc�1�&v�5����bTo�V7�M}�Q���<WH$��0�)MO���2ˎa�C��i�@ @�����]oJ�G@6�7�S���Q��)HvZN�GҦ/����Z��q�⣭O'>��,���{fJV��e���iXQ��Q���f^�h�*P�&�ʔf�%���Ew�y Eew��h�	�ؔ{��i��VK:"a7�.`�B=fpcN���i-�*'S�����Ӣ1���\����Yed\�P�'��<�"���k|��葼伐A�B�\*��Y������鬕^[�+�����K���h�5�$��9��(x%����`OQ��*A�L.�I(7U�RC���ͨ��m�|�~Pdߤ{b���`� ��"�t��r�~��8� z$eK��R݅]@�x�K�@���)��	������ɰ��VxGCP3m�ʹ����̍�j�Vl��|�c�W=&U&-����Mb�eG.`�EY����T$4����R���۱���7���_�-r~}t���:�hUa�j�K�{��3үX!UE�0�^���u���]��r� >E��~��P��0C���a��f����5��]�����i���K�����C�����(g��ܕ�y�{i=�@�;��[}��á��!g�1�u�(Io	�>?f�e�����?$:/�,3(er�(R���p[��+ �%vv8��	t��s ��~5����c'�o���@r�x�%ŁL�ϼ��p�&�f�^��]�M���e��d��ɕ1����<yҟšZ2FzC@`��TZP�]'�9"P@d�������"k� B����I���M�=��pn B�A���~�<f�m�G��{u;0���LܰD}������+��ɖ�-�Z?}�4e��:Ô3����J��1?�a���իtqw���p�+�k�8�R�z�o�KIʆ@9R�"6_v/ ��0�|[Ŭ�ʾ .��]���s�/A��7�H�o{~ΐy�2�|�.�i �l�
e5)Z��Θ��6�j�!U��,�*t({�D3N�/v�C�]�Xv?�V`� ������q�������`�jlQ<�SB���ayV3�c���bP N��DS	���Ad��4�܏8����5"��S��"��s@n٣�)�/��	u����%3�o��Ğ\�ޙ��-�t �?i!`J�,��t
��ʨ�Mb=bF��Ŝ���u�|J!�_!v�C�K�~���[�kDw��usW�����"��ċ���mG�w� ��۴��F˩��-|���B_��A.�� =�8TP��Ҋ�w��3�Xz�Jo��!��:�_�u2W��p����O�4���B
x����G��c|��Q������sD�e�U䭑R$�'��%>]�|����j;Bs�X�궫��"�X0��v�Ӈ_����{~�3�-?��CxQ�FE��>��o|���q�ݬ{R� �Ă�$�TI�ˢ]߀���t1X�z�$�M�jVl;fN`�<��Q�<����08�8n@E5�����DBm����o�ɢP�s�#5���e1��m�%٭:y�Kդ
P�ݩ�W?[a P8P��%�>1�c�` �)��Ԁ�}�:��ta��{#��7 ڡ�oR�ղ�|�H�R�g\�B�_X� ԣ�5`R7���4+�?��o�ʸ��:W7F�v|li�	��q}Ơ��)�]+�*XO*2j+m�G�@>��F�H=���v�i�Г�$�Skn<�)^�u���i��S�8�'#�2�A��Vꥅ����L�V@��b�m�6)3j��d�_w���e=�����*\'e£��,)h=�1ۋ��Q��9+(�y�*�~�TS�ͪ��ߺ&��n	H�`�k�B��1�[�q4�r����C�s��2��σO�%'ruzB�����c��4 v����R��ZC��Y���l���);̢!�a�	c�����Uy�(+|�L����x)b}�h,2���C���\IL���[(�����z���3�q@R�;��S�2g8����tW���H�t���"���~E����Pf���s
@π7\ �"�&7�Pk��N�o&��F���x��@��}��8^Gh+��g~�%'�����O�a<��fB��*��~1ً]��m��JY=EW>��F�����ߜ����l+�:���0k�y�P���9�FL|ڸ1��.�.�N�Y�4
׉�8�:�};j1�J�ܘ��?�[;�ҭ��U�7+��/G�<�W��6�x(��ǥ����4�!�ϋ­���L�}f�-����	���<V�y+�'i����B��ih2���E��7S�g��
%4�S���04�Զ/����]�Fԡ�i��Β�ɧ��ԢK7o^�޺�7A�s�ņ�j�Y<�<�Ů3�� ��m݅�_ώ���K��Ee�"��o�m���zX���]�&�;��S͵�[�ch�Ä�s9��f����P�xY�{�I�u�g?�l4�&����)X%����6-��i� p�mWF�z�{��XU)���ouM@�p��8)��,	�4v��,���u7̵�&�&��� ���)��Ar(��(U6\�5_I��,� ��b�iԉ��psx�S�Q4X�Ӌ�A�)�xx�H���S���ҪAomI_��s���l/�oo�N�)����\Jj᦯v����E�ޞ�)N�Av(���~#y��O�ʶ;vb�u�^�W�f���ĞCG�!~�#��B<4o՚LZ���$j��loDVb���V�l;����`�3\\�i���ea���d��d�rF�^2@��xx���<^�=�h��,>�*^�&B� �60x7>`��Ӷ�A&qx�p�i�#���jt�V#N�b���H��/^u�h�ʁ���F����w�<2McO)�E��&ZoNI℠��
i`AA-�%	�p.=�'��b�a7�h�
���S?�&����:;��� 	$lw���`"�F���O)?�<��cއ^`t4�.��	>�D����oY|�M��3r��g�nɭ�g��\�/�N� tw�袱Ǯ���*cFYD�PF;��s�D�����%��U`�b"���=z��4��P��w���)I�lU�{��J[���ZN�>��\��5�F5#;(R�O��las%�N�c.@d$5'F����D�Uu���ԛgǧ	��}R�-(�6:����H�`�6D�rYU�:�htk��,�{�P�3d�`�-�ۈ"�J�%���օB=8y)�)�<T�����,(b'����{���ҍ+5���	���l�g��	��K�T���� �l0�n��V����}�ζ͘OY�G���n��:�ZT3�U��I�_�Ѓy��G�_�fC�*�J�sT�0/*#|�V�����6z\����|>s�`5��.�.����f�O�ՠ��*R��P�!�l�m��/O����
`��I�D���.F\8����uA�v"������Y�$*Rx�"�Rq9� p�g��k�"Mo���1E�~5c�l�s��-2��i26�Y���r �u���-α b�l���{�G��d�E��ʝ�γ�#[U�x�S`�D�� [�)<�vT�}{�j�������wRc�8X�l�_p6�u�/:W��|�CM��U�G��	ՆL�����iع�c�V�e�R�tS�����1��m"�ɫfT�w7]ߚM�❡�h��@<�w	Ke'��5�vC�&N`R�@l�f$.�]KFe��%�jX��;�&0���L�\G ��L�vE��Z��.�{Hk��q���v8�فh4��&%]�w,З8w�ݪj�[�sj�a�Ytl�5&YY��8o?7���d^�.f��g�&3�$H�RQQc����������ܢB�#�P���bL�� |�5]�V��Ϩ��
�C�x����9j^4��cLM��ȋV�9I��g�q]�K)��Iu�w�4^w6���F+j��f�����*X{L>E�DY��N%5���Z�V���B�8��=�vJ�[���-���S�T~�N�[��3;�+[���`S(sC�j�'1���QLKzw�f��"�����a%�W^��#M�Ǿ�S��mH��,]��~���>�;a�1�q�o�	��D�F8)�%+H)�|g��* �A~�l �6��а�g��tn.U{釴, .�0�j
��@�U�K�ɂ�D�w+�.��	ݺ�����o��{^!4�O��Gފʰ�@RݭĻ8C(��N�����L�ʚU
�J�)\�q�9)d*z������p��
X�<�2z[�s@z�U�Ob���Gf�Q��O�ᳬ����j@:�wn��﯈.�͒ݏ/�ͷ�*�ڠZ��y�T��ޤ0�/���%�!d�Ν�7�tZ؀{@�Bi[bUP���o�������  ;��l\���W�
�ïj�ɍ�f�剟9��G��PB��>�:@5Ǒޚ+���@���0�).o��-Pm��ֱc|���.�1��312~��o�z  窂S�d�oT�I�J]�Fn}Eu��U5���qvwj?��9Q`&��1���������%��ɭ+��P��<�'�<��
$�0�{��_�KW�ք3�|s��F�T�W�ݐl�d�n/
���~<K��!���V�N!�YH'���Z3�e/��PiY��U�� ^�����!�r8��w#�c�(x���|=D�h���iJ��^��м*m�qC�Z�e��[���o�N��k��d���^]�d�c�����8�ӌq�P�C���r���}��gV#ecAד��V�?�{S�e�+�yo�Y���y<�j_�%��y��#�Pޘ�[}�
�Ƌ���-*�+����)�s�׿�H���Î����UAc�3�T`���X4/���zH��+?AW���� �0�
jDI�&�
����\
�!����߹�B1�{��0t8`n~�i<g�(��U�n%����3�� `>^�4��]>'� :s1PU$�ҫc�qb����F�)�vm1�{ ���U�t6;�h��D�8(� X6�Y���#{;�l�a�L<� t�2S~�M#�@R$�*�S��[��+%ܷ����r�{QI�FS�� h�H��j��/T�yQk������]����!�~��-O�(��a�)�,����&�B�b@:J�u�#>�-�K�������uۥ:��l��M5�:�W����f0%Әf�����=w�$�� #�#���V/��263�~ �����6Q�N��Y����� e���Es�b�Z�0���EXVUѣ���wv>s 8<�Z�N6	E�n��7�]�Tj6rO\�.�lP��s7��׼����K�Wb'�sa�sX��@�W7Uw P�Ve�W\�w�=G��(�x ��c\�d��:���Km����;[16��y�4��8}����G�Sk:�zk�v�6�����C�ĩ��9�@��\p"�1Dс�`�;�|����-&[۞�[...{�
@�L������gU������ ��<�Tle�Q�|:~�>�t��?g1>?B�j�L\��e��sK�1���\�S�G��������I1w���G��.���I�YkP�5�P0l�?B��9��Hki�h Ӹ�TT�o�hXJ�zH&���#���a7ŉp�n�s0�x��0��e�����-y�b@��e�
�sV���]to�}�}8\��+r"Ǐ��>�ip�&�꛺��V�
�F0�&�����E��A+�_
�`d��(��[����Q%�u؞k�A�&"�e�4]:���pW�i�x���y��Q s9c�U�@pU0$�����%=�9P�X���
�"C
�D!�����qd�>k�$�i�Ѱϻ[�b4=�˸��<�:s%�fe �vo/-��cI���kfrS���1�N?�$ͫ��[�[�Z��QJ@Q�E���w3֍8(��~�FlV
�ɮ��b�򶑜X�q�U�%��K������ɰ�(-,A�� 5h��(NʢoQ��p��{��p���+��Rp]h:��.����Hl�b��N�~������ӹǬ={`�Q��ZJ�?E�X�6�hB�)7�3�cb���= F欇
��~�9=���KhU�k�(6��Ch1�w��M� �ǀd뛏 �:�
�|�2|q~�^Q����"���6�ulK��Xа��DZ��RBjP��Gو)U��'������p�(AL�"R�S}������m)`{ NP�0���|{��B����Q>�=��ߴ9r�o5�~gx.H�)�S�T,Y�����?0l�X�{�} ���wh�ʄ���n��ą9 G��=xC8��Sv�p[����v��1c�w�_��.�^�4���M���P��z��T�'e�'��g(���x�x��@��~���V'��q��3��K���,rAu@Ej�2���]����{s��3>���anѴ��"�p��k%�A�R�&���p�?��~��� �T�q�Ƿ}v�c��m*Zb�E|��d��*���8.���׻�Ыr���i[U;���347Qv�|V�Y��B[������dG���\q��pVfNy��R8����C�ț;�ߙ�-ٵw$�.�x��F�I��M.��Q^����v�J��n����Q��\��n�;#s�6Nɳ��b���ٍ��(��i'�{p˙)�t/����Aq�e�6�!�M�b8�0 �.nSݛ�H�N�ewl�Ǟ��s;���(��� ����g�U�&�6���H����6�`�k`A;Ŗ�.�=��na��*c�T��9��V%�������Ұ�g����"�d���b4h�y�ة�M�9z�Y �9��|A�| I���G@�����:,wˠ~cCg��ޯI��=��o�NU��Ud�������>Cy�kFݸT���4�?��F[��qÅ+��� 8�gv*ix4�n��s��(�wX)G�^\��-��Mu�S�0��4ai��A��r�86�^t��v����;$�	�Ir&�����6=sH�+���4 ;�c�:z�)XRhg����`}��PR���1e��gފ'���;���h> ۘ�}��af��Ј��6�U.UC���*I�yJ
"���<���2_�G�q]FH�28BP��^�T���i��Q����ʒb�]G�-A���\�;���]0�� �A 6�����!�ۅv�JZjrt���*�kJT�4��Zu�Gʴy#۸�%����"-�����NW��*~heh�i*�?~��q��6�N)u��Q�$�u����׿u�*%��j�J��a7��X#�����i�M8)��T�.K����n�u1�gƟ��VAQF���� ��8Zp�{�h�'Z/��C��������{����q�����P@f�Y�1SVÚa��L:��ss��<��VP.z�X�^�x�?k�p�&m9�4#�'�M�P�"	��D�SMK�[��J�2���g�-�(��3:���y^��O���\G������w������������y��c��Q�����o*+|��.�t�3�e��i��6&�q�'��Q�N��c��:�`̵�X��#�����.ٟ�g��1~\#��@��@�$,ä�w����=��^��.�<��ɕ#)��W���с�S�/����}s�/,s)�D[c�dM�<��W����P��ӯ�������Kk������V��٦���y�{i�x�[��m$�A�b�@�G��<&^�e�1�ˆ����J@�%	X�/»�\���!��d{��=�v^m��c�j��/L'�j��Ώy�k[z�~��Y�_/�4B+n��e�u��Ҽ�W�ƷL3�9%��/V�2k�#)^���}lr��4�c~�z�fH�֌��ˊ�I��\�#��B�ܿ.�����������.�gB�留��@l ��L���P���=�R"�;���ww��4җ��
�~�#�]���~�̭߉g��ݪ���0��)AA�� ��'���^��BAb6��D:�����n&�l�^6G�6}�v�_~��E��@M�psX۵�W�a���8��ߝ��c��q"M��H{x
l�]|�v��f0��k�(w��IzV�踏:�<�\#%����:����x+h��jC�"C���hd:   r�yU��4�.D��K�W�n�U������W��g?�k �
�w �GĨL��&�Z
��_\d��qg�͙5�ʡ&mr�����ҏ�)1��œq��푇� V(�c����5%�1����972r�+���(���=�kQ&h�"=���ߝ׋���XK����%�o ����s�bM�ܤ����,R�f�����������L����T��+�f����u�?9�(/�-����?�f��?^Ky�M�;"q=A߈����t��2p(���'���7�qu����~*��x��I6r�(�fF�4�-��9A��y6���~o�9R��Q��<��n��n+<��6�%�t�}�F���A�I��
h������7����������P��i���TR%^�E񛰺whWW	��T;���_9!Z+gr�vs#FEV���m�jF4�� Q�&D�D�F�Z*�I��^d���#�i�	�C�\���Y��͜���&��qIȃ��#ٕ(>���қ=p{C�~1����[�қ����Z�+}[����M�ʇ�磺��xbr�Q�$�PWۉ���]{/$��_�<u�X�a��%��|���2����������Zv�Gy����ZW����.ap<��o�:�U�4�Ϗ�P�UT�a�:��T{fh�#A�w}
%
���P?m��my��7�Ct�X7zv�!�nb����m�@r�=��a�����݃����_+29�5��+��*����;m3v��k�\қ��=?>��/=j��T���5B$|	K�8ف��X<��M�hJo�H�7m��=Z����T�������h����ު��h���9lw�=.��@�3��?�����D�z�:Z�}�tݧ���@5��eN������^䋴�3��ہr`��yF�5%��ٲ>��7%&��$x��M�6'�lHz�h�{�n�ɽHUe�y�>���4�����"��g�*�����׈��!%.~� �}~��d$xL�>��,u�n���)y��f*�#��Zp������~d��J�>&��7�lMt&
;M����7�Tۼ[�����ť��4�@��Y>�`Q�/��/��#�-�n�}׳.Y��)z�E���qj��N�9��.��ؖQ���}7�m*;��Y h��;Q/��m{K�l�g�����޳R���c�	�d�F���d��I-%�����W�6|���-���M�90���S|k����S���g)��;�c�o�!Cb�П����!���E�$���=�f_�?���		�<w'$���7Iț��]ܮ�i6a�i<�Z=wky�6��x��BW<�%<z�����}�pe��� Pn��C�z,z��)o�<������+�����dc:�aj�K�AW���C����N���Q�g�mc`���,����G5�
:MO^G%'�)��F?Pt�?�'�����@|M��[�W�ժ��$Y����#�R-���Y�m��02}����S8�m��5��s�r�J��K"I� {���Ǆ�S�[�Z5�����a��%�[+��3a��lɿrT���c	�F�d�ΤU�#M�<�����n�����_-�� �b��HDTP���W���mJ�tkV��Z66:�B��\խ#
,E�Q�p4�y�i��x��L�Q&Q����Do�!z���~�E���+�D�Wv3�yϧ�N1�)�W)�x���Щ�)��T��,�*R��"e���γE�=�>-Ւ{��p�; �=x14Q�n���lqY�N]kF1
^�w {�R�M�'<&�}O�t��bF�M�l�W0D�(�]�`�j�����H�� �N�%:��
�19H6]՟�@c�b������H?�h��EW�|�"w[O+��=@ Q22�F�����k'�q��:_�(Ķ����7M1�y�n�_��:{���L��d��/�R��O��ف�Z���{��^XU-B�a;�'l
���9���A�4R>`@{+깞��q.�'�w��{e�\ؼp�t�+7C䉃���چL�C_���_�J5�U�_�pZ�_�����$�	���8�o��R�@�,8��6��hU�Wn+�T�W�J��0�[�tɵ�Fԧ�>H��!�(^� t�7d�@ �(B]��A]J�^����O\����w���`E��d�\��pN,aN$���M�{R|���Q��[	BS��f���g2�7Qj�IǝfZҔ��� Q�D׋Az�)"���:EC���E�̬��m=�8{��Kc���hg獑�6�꥚�A]	D��3���X����@������88�m�J�A��!�����%��~�1���R�y ��)"��l\l��
�f��g�b[l��mZ�[�)�o1,�Ծ��/�k�83?h������д�Т��+���X��#�g�d�&Ф4'�w������J�H�5)˹�&�����:�B#�n1D��G���r8���i��)� �=���>^	��e����  �0�ԟ����L.�Iq�%ʡ�[����6.ǣ�~6��Nm'+�*	ß��;�
���:��9Kڌ���)<����3��u]�v�କ��'l�%�_t��H�}.�)�Ю⹅�8C���8X񒟎�u�w^��mf��]R�e�ӉB�/��r/�$��.f�l����1L�ic�2�P����
��t�T�er�IrE>:�RT=�eՓvc"��?�Դ���Y���F��F�3>�}|�&2��,�PنiR5(|X��Ixtv��0���mJ?������w�[�q�60}�XI����n�ަl%�<��s�?
 ט"��|v�06�g�B��l� ������i� �Ɋ�#����wk��=�dh|)&���*o �e���Aǐ��M��MY=|�0���>O�L��4�+�b�bu�ew�a�7+p�=��;Zy\Im��,��G�4;AkNO^�fSb�[�ߺ�p��I��^T�Jn|%}\@9igڜp�����֫g�~��Z�Np@�ui�jA'lv��-��s���2�,������)1��h[��5f=Ő��j{��joψ�������hl]������˄�����WwLSk�ԝ�v�x�K��n;}�Y�8>?�h�ȫ�^ ��������6��az��(���&���S�S7��g�Ğe�%O'�3����PEA��m35ĩAR�����{
�T���x�'�@���cSt���sZ��3�@��V��N���kK����ӆ���Z�<Nq|2�N��6����z�� ���	$���S��OW������Rl^]��{�3M�w@:	�y!G�N��5<��Dn�Wr<�U���Ax�Qd$��0�ڰ�P�Ʒ<���{���������1�b��&6Ʌ2��6��v���P �z�ʷ���ui���	 J8��w�э`:�e4���S�]�,Z�Y��#�</���Gh?"o�(Ca�v<G���Q8�C@���@�}GAw6��un{ސ�kCxsH�P~���_��I�.P1��*;,Ӡ����ZB��1R G1j\ٔ`�}ԁ� �����m�Ȍ�;{l����ߵ��y:a=4��FO�Z�J������FrLE$�/C<(9E/�t`>2N�Sn3����6/Ja�N�λ�@����y��r*ZkrN,PH�0b��ĽUKM�j�{�fo�����*F�x)�w�m!
����X���r�p#�@�
�&:B�/��s�ZGP�.N��r�X`�����~7j���-)�\1&@4��I��mE��3������
�����wq	w󒞮�5��)�1Դ���]w����N���!�t�5$˄� ����Q����ˀ�x����E�N�r�*)��o����q�L}�p�p
@�����7�eO�� LC!�48�`�< �N�!�Ȯk��ϫp��������Ք׌�r����bb���0dlZ4㠄����r:l�^ Ud��u����c�Jb3K�G�r��Oߠ���uw&��60�y�J"�B&8����\��ү�g�,ݜ,}s=�A�ͪ�w	n�&`�0@9l��g���\J�5�>���Į^���z;#K9�W��H�^$N��DEV6R���D���&#�@<�����ڣG�	�e�1kn�b�_�D%��F+L��q����X�x<��?-�7v$�ί��vX�qS>}�|����?��T�e���~Au:�pХ�a%�现��s�XǠ�k�q_y����q�J���$����\��u+P��u�x��b�U_�?<�ͷ��P(bmg��k��E�蕺t�g�{)o&���7<�W&䴑��a������a�@�q�5�Tl=���������6�e%�+1��w�;�Fn�$�'��e���IZO(��2�q�W�d+&�h�A�R]��:�Ll��w��r��t��8[x��a�O4�HEK�`�D�HV�Dd��Ü#���CDgx�-�R[Y�ҫT�͉��/�uC�d}�Y�{��v�:��_=����»Ʀ9}����Y�x��Wn�H>�`�2�V��k�~|���$��W<�3>����Rm|�Ia�}�f����09������Ry��!N����n;�� ���%���0��#��5@��:!l8�}*���մ�$����Zi8L�Jx�|�XR�="�����^V�J$����Ǚ��!'Q�Dћ��2&�^V��3E��P�^ut0����w���&�ꟳ���o����7�{���6�v�����ܾ�Z�IJ�`ܷ˓KK�㷝���P�-��������/V"�=�<>m�n�|R��%���ڦˍ������[���8�~�~,�(�x�����\�y������}��6��h�"r�F�h����լ�[�	��AK"zB	7��_���]��x.v��q_H%�����Ve�>,�%�/ ��O^�2��699	'kk�gP�,���_���낿��{��O��է��Wk�X�~*Qw`�n(���xٝ�(�`=��_�<^�)��+?
铈v��Jz6i��[�H���v���Nq4�ޝ�X@��;*��M��Q-z�޺,���Eo���d�?�$Iſ`bd{�Y���'��g`�]	���,pӠުVz+>ش�gv<r_�(к�r����H�c��1/M��&��kc1z����lI��d��$���t�~	�M�r��ƣ����T~��6�L�}�(>��q;+~Y������-&`�k9Z�;�Jjn��r�k-I!����7a��;��`�q��gV�^��		�~ �W%}��7s�\�^�4"^�P!Xp�ŉS֧`a�)���q�.1!$]��b*D��C:�~k���EU�h�&�8��m�������K>��s��'DQ�m����0/W���|�^�(T���B(�����)����_��"4�����}|ȣw��HWb�u��b�%Pgљ�Tj�m0��������)݃]_�5��'x�Q���P��J��J����B��ܽ�fo>Ҷy3�ԮQSE�t��"�<�|�J-���n��M-�ih�a�H��-�~o�Q��א�wW���Y�l��2v�)����Y�ˢ�a[�������A��[��v����8��>����~�A2k*���Ro뙄��ڝ�^�X~���t����f����gn��@�����[sР	�?0_:��}�?�s���r���O@�>4�����{<[�ܵ,��581�8�<|����� ���ʎ�B���0Y�;�!��S3C{o���[SFʌ5�6�d$�����om-o6�lX(�Ѝ��|��L�����χ�~įZ<�[s�����;n�F���Ӷq� ����:�m����B�T�: ��<B���+�͍YW�  ����\��5P ͧ|1A8��+���QE���ߋ����P��+	�e�8��oW �b��%��!�V�����j�*-�Z���*�c�N0X@{u���-�R��M��.�}-���V��z��`����a>n[f�~ޡF7�e�i{�a�h�2�����B�N�Е���5����c���y7;��q�9��Ԃ�G�7!\O�
:O*yZ���<��Q
�r���a�d�h1׍�Df�d�V�g�Lo�_s������_��,g�HY�ϒ3�z�:SBxʩ���X1ئl>QϮ'�|��oX�̥>����iW*�K�P8���f�Mz�/+;�/��#)����]7ʥ��D7�9+�f�9x���m_Θ.K���_ٯ�΂����y~�w7���犞�YV�[�9i6���`׍�#�O�wqQ���s�up��[^G�9�	�;�"g�5�6��4@�=D��6�P��j�!�����t@����}�A�\�\�*����Gw�R�O��Y�s���S��hau�&P-6�E�jOog�c����-B��C�(bu���è ��;��{l�i��P]����__P�v���_�nctr�6�OI�����'a�M8}ڽ��y��-�$L&�ڜ����Y����.��X3;�p��Do��o{*v���!��)%�>�;n��ӂX�%Q���;<��H{��T����=�a.ǒ��|H"���:��ݻ.?J��2��}E����f�AS�
����{I�OK�2�=�wOZ��֮Mul���:xk����z{v,]r鞠�4<��0���&�Ojaiσw�z��XG��T��
9��J�ڹ�9Y�xQ�ǯ_n��k���3z�;V8�1S1$��c?΀������XY���DT�2_���\E��aw%-|y�((���9V`s7���i>�����	k�ZB�ʶ��n��J��E��J�b+�ʺX�2*��'�h�{�X��.Hfbb�&1|2��J�Z�C���qǐ,�Һ�(Y�������ֻ��۪]م����5"y^P��ܰc��l�L�<#ʨt`�3��?Q{�y���/C�m���.$�%o���fW��1�L��P+���W����߼�����pz��9��	;?�k}<dٮ�y�{!0��e6�d�M��Yxv���&�Ѝ֧?�bA8���ξ'%�o"j�����h��Z>�������"Yd�uɤ����9#v��q�`�K�������ܝh`��������P1%�o�9���dd�r�������U���>wMTD�h7�${u����F�K�Ŝ��#�No��I��5y��n��Lϟo�>�T�sd1��~���̃�9���)�wWhsP��fJ��π��\��ؖ�)p�h�>��*إ팲�ٟX���X9��10&KOÑ��u�;�./�E������������Z�O�Yʵv����R���{ۆc�k󢹶"��CNB	3 �m.���/�%FeW����_���lzk�� ��ɷ���ѿ\z�Z�z����ZC!�y�� 
�}>S�;0cg��,�%��������x�f��ȉk ��>�o"�(S�&�@��>���΀���}k8�
�D9]�G�_/�`S���������~a�)^!��iq�.,���vBn6�32���1^J^[?���دqq����0<�t�σ]$M������ 0%��B��'�g�4��X�r����Qi�\z:�3��>�:S�rf<�B*q�ء���	��
rog��x��4{���	�;^�@rھ��k���[QG�,g�>����"�J��ij/7WH�]G�D����5?�K���i�x
sz�d��!��I\ps:��\�67����be�͍�.��L��b��%q�g�^�����ޤ
Ck5q���o��">@=Aɭ����e�1�Ř��3��ԉ2�����B���azJ����/�o�gh?-_	���=�$BI���.�����v�~_���3��\���Ə1>6��o7)d�a�����_��� +������x+�?V�/N��}Wl�����9�'J[˞jM��U]���j�j&l�?��ߦ��$?˳y�IM�l��A������#3�4"�%�V�Ь���
�}�ߧ�]O?��H�pnI<�ы�e�����?���U���#�}���r��v�e_'Q�;�#1Э����+�Am�o>�/����O&ڐ#�$E�C�����ݔ�O�B~:���7]�\JD��q�c�E��gY�\q?�>`�L?unMj��p�RJ&p��H�m��:���6��O.��Lf�ç"��^�,qo�h�L +Q�e�ݨ��,�I�2ɛ�;�C�YXb�0�=����S�8Wµ�Y�r�}��P��= 5��%�%dGv{T��C��J�c�jdn0<OM�Q����Y����w�S�ˈ����	/��}�k�c���g�k������=g �K�^�PKD��u���Jk��n{� 0Y����b��׵e"!�=�z��l�o7�#�!��E2{	�^m�}�J��Gu���ҭ}��V+�4>"� �
2��;�I\�s�����'�v�*z�,�O�1��]C���v7�~?z�.� ؾ���ω	�]?n�{裏˒-��/Zy��PepQ�M�R��\D�Į�^*g��r��7~D<$�H��>��{���I����0���x��'����o���[8W*�92�?*�:.��k�n���������N�f��i�;����F�T�������O<sf���Yϳ��*{YI�$*� ��z�&��O�*g�=�Ki�Zm���ك޿�*��pAK.�@�2<,�~D�s��w�_�G�{������%����;%;��*����@�@᱓��Bu�C���"jB�ʇB�Ǘ�FO�C�ͦ!D��Vo�8�2m��wъ���U���`�z*��#h�>k���4�,��nt���lO���|U�G#�~�`a���xI�r,|L�$Zڛ�G�9���%x�w/�j3&}��2ނ�h�S�yi��:T{���/��C��ĨDil��w�޴P��$��=|��̖=����Zw��7:�>�g0~��\:r�8#,t��hx]d{p|��c{�JX㢅�I�)�8�ȿ��h�w�%w,EY�҂����7D��ɭ����>��k����2�Z%����i5B�V�5p<�K)/��H�r�yuy��{p�|uV���}��r����)��[kD�/&������`�(���ThWDg�Q�!5���ϗ^�.Ds"ZГ	s5s���|��!y.�֩��a�`$����׍�T�ter��p�@�Q4�A`Fϋ9������y�f�h�Q'��(b�>��ĵNl n�G֚S�
�I��4�\L3�-S��O���f��lS賴|��5z�oL��ڹ��;�'�b P��
<�WK;�B�K� ��������Q�U%��Ǽ���,jz�M����+ <P��`1~*z3���~I;*�����,�3\��"׷(�t��1O�G[509A��]A(^	3�Yi$�d��-�Â��;�]��N@~[8;�W���jX��-�{�NŲ��{����(��?Kb�Y1�Y�ՕOi3�C0��j�o��X�5w��ϟ�O/���B��n��;:��({zY����	��/h��>{�@�a�GS"%�/Y��*����:�%�b�*~���J��џJ?P�;5�,lY�?�j�A:�R�#һY�/?�cW����Ǟ�)[�y�
<6�?��o�5����
�{������H��s��nh3=G�-�F����)���n��;���_��jSʎy�_ȷ  �ΰb>�LU -��M�s�l�"R�ă�;ڥ��/���w}]fXk<!2#p����#�mqδ����E���3�G�ivX�B�;�A9���Z����f��xv��M�T��]H-~�U�kZN�a'��b-�����-�]�������������aț13�xam��G�K�
g�{����c��m�j�-B鄬�����Fs�Q0��h�U�n��wc�!�0��;*]K���E�Nt���g�d't�T�j���'L[�� �ɿ� �2.�ߵ�j�(ǌ<��AZ���������JZ�b��Z���m��=���Yo�#
7��*q;%���y��Ij ����^-w�UO0��,��V���F����Y�m��s�K��yy�D�y~�M��[���T�=!�`��E�Ƕ
����_��;���r���O�ϟ�y�w0Z�Pc�Fh�5�rsh5C�y��j������j�pې�3�HF�0�(��n���Z8����8�����/��0�K�~0��%m;���r��ƶ�ܻ�J��y�C��õ@p(ll�m��z��v�H��-ܙ;���Z��E�:���TL�v�9ò+W��e�G�\�&(߲I>�FI�,�3�i��W��M�� �Fg��k؅�}�u�ZNz7�{IN3:��i�ń������e�(՞
IQ�`�{g��++��x4U�{z�C�M;�u���]�^�7�t4)�T�������FdX��-����Z�aҙ�L�fW ����@�3޳I�%�_ˈ���a'���.��+C{Ѓ��y�a�8V�8�R�1�kU�1�2rAٓ��I4���xSP�uqf���p<��h����:�i���N
K;�z%�t%�ÈKh���m����3&AF=�ύ����|���Z2!<=��w5X���I�-�(���B�u� 
QA}v�y�'�3Ib�8%��:��S�����;��{AGJyY1XE�XG�� �/rn;	l6��MX}��S�Ki!f���=8�t�'d�:[���#�v6ƚ�����\�Q�B'0ʊ�S�*��]��ۭ�!b�E��k5���/;E�u�4hح�7��G�:��<�Y9}k�/���-v�w͸�� ]�Yu�_�G�
	�k�q�Z�^��u��h?}�"�ת�ޛ�����5fmX� k{3!�$��|ܾ�Vk�OL�QÅ�׭�tZ
�v�6�
����EEj��}��?�nt��*m	�}��G�yk�d�ff��`�9�r;�o��2�,�-��ܱ��tF�a�f�`�`��Of�wCP��]?ZU�rD��G*��~,'�D���f��{Z]P� ��@��^ՇpvQ9n �!}��z4Х{'��D���4̸�շ0�26��ܭ�'�6��k$�&�%�]烇��^.�j�cP~�Dշ���]�T}<��'|�����ź��'NK8HU)��ufO�#t ���KpZ:4�p'�I�I�jU��<p觽�&G���LP�d�"��猒�����ߙ9 @�=47V��u��k��%U�Xh���A���"_�h���˙U��N���F��ݴ�;�]de� ����f���F��#�z?3Ge���q.&��8�6�Vbq8
�!�j7v|�ub=������ئ?�>�h������%��w�5F�� ��J�JB��RF|��X�'�����6��_,��Cv� "R0{��.�T�nQw�{��h�}i�򭖞8?Nٽ?[n,�ć�(kDʀ��A��}���Գ�S� �ȕ�&�
�'�������Gnn��u��ă�G|3Ih,��Q$l3K��r:x�O���^�������t�*�eg�_\�I�#fj��?jXO�5����l*T����z֬˶�uo͍�h8-�q�Lbge\V}xt�Ĳ�@͍u��3��ʆ}���	�����_5��?�4�onԠ��;�?�N������T�%����1��2P��)�������]vC0N��PFW����������x��������4:���������!���q����� �dJ�=غ|�s�Q�u�4�d��C�X�2c�p���{m���l)��XI��ˊ %�&��8h3���楣�58QNi\'���������@3�z�]��t8�1��C�Mf�W>���������O�np{��a�Kb�1�,H�QR��kJ�Qإ��(r3I,-U�Y�s�pZ���M��Є4�	b�sr�:�B��Ч+��蒅P���>'�^�����7+)�_++�qU?��z9 ���.�~k8���>3|�ʸ�������5�4���[ٝ�B) u���tge
�b���h\��R �ȫ�wg��x&QӨV8��dN�s]|Nt���l�D���=��g�a��,
w�f����o 3�<n�{� ���M��5����\���=��*И�fv�KO�'��fa�7U�l4��t݅$�)�����bh���WhgH�G@��4V��|/:�H�<A!�҇_l&�'�]
��/|R�����s�M����uy���g��Wy�ȣ)m�v���z3h2)��45�)?Ί'P�h��7D����@}���@� �[f����{56�#ͦWg1~B�I�"��<��E:=p2k9�R��Ѹ�Cnz��f�QU�hT����}G���#��V	|M�2qa$�XJ˝,;U����f�6ۇ�P��M_�&VxqTe�C4��p�����&9�m�~���v�t�g����߼4m ����T�u1=����.��1�V��O0��@Q[h����F�}��_3�0!<[�ǣ�-�'��{S�&uԂ���J�� l�5��U$Ф|�s@x�L RBj7?�u|�z�,���l(@H���T�����07����.Xʄ}UD�U���_+�9�Ä�6�d�2�l�VV����r��#X��ߠr�\��Q#�R0E�fX��gu� 0�������e�>t�d�
�h��?���44m����6�M�D
�QF	���)	�i{��������8�$��?�����M��UGY��B��k)F ��jj"��u���\nI�V]��Ȼ�\�o��Z���3���EkFw��q|��®���{6��T#�E����L�]#��h����.��!�h;��û��*�>��|m�
��j����3}%v4��ӳ:��C�R�P�6�t8�x�;;�>%|��P>v>d(�h��v'��������t�jZ��F���_�6��<��X� ����,x�X6�@}���<�~��!�o���o�y����&��%iQ5f��3I�ͻƫ����L�>�7�(:LA��(�qw��r�/�u+��x����;�>]<������t��D�����uN�p����!u���E
�������������!O�eC��� ��J���$]-����$�W��y��O7��zc�=0��f,�5���D��t>rbZ��Vj#�'��l��@���"�\@E�Cv��2���u;j+<E�9E��fm,ַ�o ��ο��q�6�RY��6$
`Ҧ�	�$�;���t�,�^=��z��O�7^��י����*����L=�oX��]U�P{_P�id�>��o��r*d;*��t/�2[�6�7�ß�.3ᯏ�0�5�����������T�[T�E��n���Qa%R���Y��Uu�Yl�o(��=���*l4�zk
"�Bթ�����������"G촭F~r��{/�S:ܗ�[�lh/Kh��7�[���~͈�aes���(=�v�\ſS��^�Nz��.~:�Rk�q�V���?��E��7��t��~:3͌��i��BQ=c�K�;�jc��P��_������ǌ�a�>m�-��?˳6h�W��������HK���oG����Ǆ�ֿ��(o�t��A�q��ʹ=�6M4�'7�c�O��*�s����̷tk%�X)�d=4�  PT��	����Mzk�F;��?�f�T�p�&��t���x�:�?�9���9����3+��D��f��(��H��(?g�+�
 �򇢄�����w�,�̌.�����<<I!N<���B ����/��C�:�W��S�l��	�-�ߓ�����p�d�(�Y����N�'��$l��lf�V}A	,��ݴȗ��L:d�s{7m���Q�/���L������e���^�|)�0Ш{�,|~�OQ E3���Ϸ�U1��n�{�5��|(��u�FGk6~.�{�v��{0��t�z�Uږ�y�k�Z=f*t���UD0�1'z�J��~�����[�3R�xk����Q
���2�2\�6@!�j�͕�lr>o_�"�v�H��T�9��XO[!�?�������0R���a/T�T��d	:|�vҠ��*���2���s�"�� O	�"T� �r?���^FيT�N���r�9*&�L�,x�s�z�%xi�y�5Y��h��qE_����v����Vae�{�x9���"�#b�{si|�?`���aѲ]Z��'I�N��n6Rz��yk��z�,�C��m�QU��3P?vH����#�X�j��ܽ��F�5�!C��j�d��	=˵�Syot��v����d�Ǻ��w��^:6z� jGֱJ��$tmuR ���Y���%6�?UO0K4��JGHB�1s[#��O�Jln���~w�3��?i8��[Q���!� y�u��z���/.�"���&9X���Շ�{砏c�����V_s8�5S�o$���FhP�/���Xŏg�����4�P�6����'"�{��_��m:��k�7��s$�D	�����%�iO����by�/��=���>��|	�D�^9�we��w>�fD�n|�X��N����Q\�$�%r��/h�d�c*2! +EB�<;<�>й���Ul�ނOw��} �.��n�y�FС��#���H��/ן�C!I�3��w߶���g6lG�(�~�#T`�ع�Ŕ��L�+��Z��K�4���� ��m��5?��( ������t�Y̮ƾ�����^�Qʘ��l��l��I�J��;�	��k��F��!+h�	b=�����*	�2}U<������Q�G��-g�����2P ��{>���pz� ;ԯ����澍�����P���Pca4Q&/����X�m���
�<K�NҜ!F�S:d�����mģu67�	xS'���l�Fe[1��O-��ՑZztk���h�L8˘l[�(�7{�p_-�}yZ�� Ľ s ��c��{<�k�9�J��e�����{q��.�;�0�s�{������� ��9uy�:�?e�=�/�������}\���
��?C��������&����������+p�&$.zi�Ysu���EW^ns � �h�.����%���s����be}!��-�~���c Yl��p�
�xܐ��d#����In9a?|s���SFR�|BM���_gW3�T��Q��/�4D��#8�FXk���]5Jţ"�������L�<��Y�N�����+C������Hõ{��c��"Ȉ��Rg#��ǝc=�h Q�3���批D2�^�e}Λ�s���E��P�O��J�z�E���U�.ms�2�����& (,�.�Z6j�)��㺋3�
^��H0��䣭��������.@׶��!	�zN��1�W�W1���C�u{�g�op�SdT�ʾ�l_R愯ow���4㰦[l(���j�e���%n���p��F���E���U�����@�:�+��ʰ�0(��� ,!�L�|�Y�&)7[
z��{�W��y�AT#r�4Z�[�(���٧�����h�E�c��.�^�ʙ:}��H�s{-�C�.���9t�-�?Gd�m=iJ��\��J����a��a�����%@��n��k��R3q�/&�V
j	�����#͌�d�I�	�\��	����Pz8��=�l�7�'�� ���5aE�ކI�\]�@�"J`l֟L�*�O,�t�(� 7ԍ��'��g 6N���5(����G���!q���[�C5�� [&���4{�����C��Q�h@�;������cr%�y���QЛ�`a�p�X�@�Ǜɝ
U�镙���5��q�F���˵#w�^��Mbg��Nf��n��#N|_�8��3���?dՕ;H���o��;��S���N����I�!S#aB���"���G�׏������,�&IW�wP���|��&U�a}}y�ߠԉ|�P������ ��������.3c�=��(���8�Z��O�o�3\ʺiD�b�W��PĊ �c|?9��������/�e�����8u�
G�yB'�Տ��)�S,���.(c?�M�Z�p ������gݣK��i�B�Oi�!��\>.�8�0��K���RZ ?23���~`)ݱ���;�LB��:�10kt�g�s���|�9��b���������oQ��	Ǉ�/ �6��8�^��n^���ᗖ����GJ���C��D3���ԁX�s��������ו]��	��;9{{}��i���2k9�A�ڹ�Ŷ��:�[_�)�S����3d^MvѮ�46���B�G=���/�e�Ԙ���tcc����j.~��	}x��#A:��d���k@���>ʐ66Ճ�'x�!V�N!폶_�^�3�������:T�m�;Z>�x�����F�u].g����x5f?1H�pN�+t,�JJC��ĕ����/�Fl���=`���㱽eo��UN�����8}��ik^J6��F��
g����m�;��=�?Ȟg�%�:������;_:�՚t���Ո��)E?B�P�K��ȓ|}'�*�$����㾕���i]%m��2��5���b�����O���c��ʯ.��c5�$q�F��Lx����*��[,����[fT4�����$��߽s:m+�bJ�.I,W"!������ŉ�W0� <�������BHRÑE��(+��f>�1��q=��O�ɺ�2N��*_�v�\с�)��ah���+�a�&� �K�U���9Ga�)W�\�?ƫZ;S�7�?9�y�c��#ַ��F� I��-���Gj � B��qaw��@�0"���{���I?�NX�g1�$I\���E��Qz��1�\����
%'��1T.]�o�G�7g�s� �X�Mw%�y.h.B�I����LT��v�����������%�ķ�W?�w�^�9K,��S<�pۺ]���'|��x�� /S`��8������O�U��f�q����� �`�%�>c"a(K��ڱ�"0cuRS��8���4u�.�$��[���q�z��|o�2��C��D\�����o����sd�%yR����6.�z�Yyp��s�?:Px�oQ��O�۽<w'= �B*��,�˟�]�/J*��oP���8�����&�1�Wj����h#��.FB�7W 7�P����=4�'!W.��M)s�^����F�t�i��S�27�|���?��?P�޼��Ժ �J��q�u��D|PN=u�s���'�e�zo��@�N'���$�qO�8Q�V0��Hx���Ga�ߺ~Z.{ﰹ�X`'�"�}��B	n�Tc�j�ۺ�C��ύ���_8�b�{� A,�v�d{�}�B�u$����P�A����i��N3\o��7�aZr�4��;�)ʇ�T�e����
�}�S5��	oG����;���s���M��{N� �����8�,&�c�1��2������̑��-��-�B5Q|�1�F$M{½��qc���~ى�1�&���� ê1(�i�I�׽�_9��锿1�籨5�w0S���xxܾ?��������:��E�	e���wa�a6�������i[6�1t��I�Lx����K�t���-��=�w �&�G3�<��ё�K$��:�]@-BAj��u=���PQV]o�Ã	�^� �@	2�WK�Kɬ�Q؄�p'�@Y�|ٲ�A� 8F����G�b��6��?L۹/�c<Q"|5���ֳ���z���� +i���jْ}ȓ���Qkf����o�q.r�ZrV�!�����b����
m4�̯A�e����o� ���}��+��#��]8ȏ�5���lw�7)�@c�
Mb/�B 3��1�1���R����7]|z�9V�0��j���z5}���0 D�� 
zgQ�P31���Lj�K6����0������R;�F���W�V�j,�����Q'��}��W��c�����K� I���'H�ʕ�Y��|�	`�EEu�8�`q�G�`2�O�N���NL�1��B�A�<;�6v"�R/�X��P���W�Hh�|���A���d�p�#g�ѕ
�����*@
3މ���t�(�� �K}����5�xPN�)'R�8Dc$�c�R�W�|�4Γ&S����>������c�XU�o�w���?�˚��ߡ��2�[�������u��@w�I���� �1�C9j��%g��ww`=��Eki����nm}�պX����k��נJ<�/Xzg,0A���RQ�pVUH�F$�K�74��\�.�� ͷp\��5���p�����e�b�0�%5�˕��������0��E��9*d6}��U��
*�Q�a�A�RAML�ef6����k)�t|�f$�p��g/�N�i��洝�h#�y"ѳ�-��'��g-x6��X�L/�5r�?9v�+9���8����&ۛ�L���-����2P�s���D��c����mŗ�d���ȇ��2�y��mG���,�gD��xPF/�x�=ypFF|6��y��$�s$L�����BF0_XR����F�y�<��?�&~�%��7j]Q�4�oW�k~�RZV�E��G����[~L�ɂ��Q꤮b�n�pf'R(���w��H�z�����p
���z�#6y����b�~�Z�Ņ�#�e6A���z�ŵk&|�!���"�2������B@��'"B��qh��	ٸ}?`�Ó�hB�Z�GF3�п���o���*D�:��Jnp�ҽc4[Ž�L�,G��ӧq\H���h%|�|�T㞴,�{�T=�1.-����o5gL�Vr�v6��c�p7���!��nNhw?��zE���$���e;m7��W(�uG z���'��}�H��䮥�X�w2��v��2��1���W�����3\eVP�n^�̓D��6�T�Lx�7��y[�FQlDq	K�I��m�@�,o��r�ց\V���|�A�lk���ύ�8']�sǑ7|�?��mx���Q�.������������Ο__�3��0Y&d��!�wN%/�i"�)��3C��u�C���.�t��$^5�S��^���o��i������+Kl���n��ay٧�<�9�U�1�����i��uȢR�A.���X}�Jܧ
q�����&ja�\م��	��j7��t%?M"�h�RZ�
�r3N0:^}���Xt0LxL&�3�F(�g+jE�2�s��I�N��Dߨ3�d�
Z6��VnR9/��'���"?-s�]��ݺm&;T��&ZV�k3Q�{Z��cq5���D���W^�4U]�y^��@!2踶`Qz�����'՜��]ƙy�����C�;��?g���¸(^���'�i�&�1	�#ʵ0=�l6>l4˖
�i�ؐ�S7�v�_s��7|J�)�
�RY\TŰ�'�DK,rN���(��4.�8��'M83�0r(C�uB(��r����fXep%5Hd1�3+r@�>�� ��?�j��?)���'O6��|ص`�_��01�9>�w�����5���><�Qv��q�C�|�P�06YM\oR;J��+�����/���#��tD��v��Cz�,{���Z�L��i�m���h���sE~|\%��T%_�����o.��M<�>g@>�k�QVr�b!��ZR��T̾i{�$�G�G���/�uX'6�[?d���]�<~�}E[��0�پХ�/�9'�c'����7V�֙��.>�ʥ�ER�-@�=���������+Έ�c@��(U��̊�v�#'d��U�'.�pT/�\KY+L]Z�j���b������hIed�ܿ_4��� ���FI������5�7���Vu�:��*�3}�d��/#�}_A��8��}���
�и1����e�ФjN�e��olA�	��p��}}'Ld��Uڬr��"u!.�B���*n�NN[�4���{�x�F	�j��0�(�:|\eK"R��2#�5���MbxV����g����إ�r���M���l�����Q\w�$��R�\cZ�������|���ʚ��y���pQUæ(Y�!��������S#���3�oE�T*-k)N�ΏV�#��}�?:�W��w�@�kyZi��}܉��>Ts��&�c5�������T jΰ`ȿ򭵣�{�!��.w��n�ɫK3/��a���mlTEX<�3�V?�ų��o^'�!/�з�����+�N�o��A1��Mu{w�$%��f�\3Z_�*�Y:ОY�[�Tpp/��s3�t#l��Q�thߪ�	��c����U`�C�W��T���J�O�fp���w?1�tDS���4�r��W ���D8:��q��@S0�mC,A��س%�1R�=����w�g�;�h����5db�N�cU�/�?]�~AS�t8�f�V�ĥ�@*><�]#"~T���0�;��|��hn�J4�W�6C�Pvt�K>K�Θ5�����E���KU���{[��� ��G`��_����7�(Z"S8�*ݡ�k9-��uD
[�� ��"m?�p{�t��^ ��T�����*7O=ѮK�6���*.Һ6Ц�p��N�?!��-��U8�3��>_)����1�;k��3&/�M���Ir[��O�p�΍2+��6��a�X���7v�5�V� ��!yx��'�kc�w��n����L�Bޒ�S�O]Fjb zpμ@�C�c�)�FF1m2�]�oq���="�>
��|�d��(Y)|9��F��Q�.�4i�Js��]²���.�̅�#;>#U]p\�}�b��izd9Ê�ą��n8�G����~��=Q��,W[ꈈEr��/�x��7�-I�c~aGBܬ��@�X�1'T}?���u��K����7���Ŏa�^w'�^����YЋ���T@����ۧ
弯��Y�/�A ��F_���mh��4�Q�˒F�-�t;�|L�<���!P{�'j(P���b!� a���/k0�� Y14��bhe��]��/F���P0��Z�3Z�?��yLx����ckSw��H����Ǔ� qW
)�R�nS���h������s�8��+�e
��i�~�NRiY'	�=E�z��_�H�_J���u3\�~+����a�N3x0���z�w�)9�GN=~��j�kk!3'G�f4[�˟��p��ɠ�߀��^KfČL�񢵷��da^�X`y �� ���Q��y����c��eX�_��g�	�%� |������k�k�)��x6�Ƚ��*U{ܿ�쓑��V��%��r�7u˟+P�,66�_�kR|��ʸh��oħbI���#J2�5��C�+�̿��v2Ė����G{tt �n-3r1U���"���_OV��[g'{��7��b�)ĩ��mĐyG��x�in���7;�U�d9e��-c���Ö	c�wҿ�V�]�_R$�v|���Q���+'8%[��n>C��y
�k�{���5�<�� N�檫�~637�M�?�8=�+��:?�2��.mn�Ww�q���ml��0a�#�h���"rmv�=��s�NO�8���g��0x��5�%崭�6�3K���'w���ͯ�����s �g_�e��M��D_]�ƅ&Pӗ�����
�~��s�T(�y���BX����m�/o�]�Z�0�ȏ��C�{G�EY�<�4��FY-�*L���A�����}��2���#�`���nyq��v���
�"p�����ٯ������M0��,>��=��!�s�*7�k�ZY[-'F[s��9:{�:0C���lZ�A��䑆�^�"X�3�J���ԣL�ĭW�V�+Љ�l�had�Ɉ�9dxt=���W���dEa����9bFR���jM�H��4���ޖ9X����'��a������
�e�����[m���~6��4׉��V��z�%C����*�܄<�J��̀�p�8�y�-����m��Ķ	��@�t�	�[蹠.'���B�GK���f�+\���E�MUa�}�V���Rdk
��WTC�.��V9����*�Vf�v��9��7"c�-�y+��aA}kÎ����6_���ʕ��{�X�׸���~��y��L��F����P#�C�`��p��	Z�)9��xk�-2�G��r�o�M�m�k x�*r��=�i(o�"�;L6ف����D�H�����^��"��(O�?��!�ʪ��� | e���#F�i٢�*�|ޘ �7_�o�ݔ{oZ���9����{�qH\�(�>�!y%���hG{�w����l*������X�?N��.��ς<[���[�1c^~i�F�V�y��u:�@�b]�.L�A�IFx�u�s�����	+�Bi!�O6�\��?��� �g�⫰�ckk�~R<���&����K>�C�@Y6��)��>�ݖPu��zE�pf�3��}q6�S����0� �ӷ�t
Xb��,)�H�o*K�n�t%�{��
[��ū�˕jo�a�pT Zh}���M���qǹ��V���5��� K��3�Y~Ќ[΅h�1�fu]E�z�
�>��$)�M��[��Y�����v�(�0,��!*I~�E��{���$*����;s�
�1�=������Bp0#����ɁL�v��S��q�4%%�T�~;�D#E��j��"H�·�۞O�-
K�ad�ٕ��}@%����f�$�zk�����5�/��7#G}i�]ƣz[���D`M����]�E����q��V�i>��	����HÑ���Y@�F��D{;�8A��Ө�����!μ}\����I��%l[L.�R"s?� ���%K?�S���V����G��/�	b����"��}�9���5;��$��Ra��YI6��#���:P��ɮp�^��II�A�@(�y�y�P��V%�阢ITpc�
U������&��]��B{g��#�S����f���``���M��[��Ӏۆ�O��k��$/�-�:e��u%�%�D�{����jQ��~)6�p,,j���ON��:!K��54)6#��,{��	���b���#��]�(��t�B���Dc�o�H��d�?+�Eڊ?�U���lS
�,�H�y�+���CgpDʎ�L����,��K�x�.,�N)��߻ [��j1�٭��?� �0�=�%RC���a�ɊXP۷��3C���r$��H�*����Z qmo�ʚL�2eϽ�)�<Ľ.�N��.H�b),��1� ���l�-�J�RP�3k�D�QO���"�E���È-C������A�>nK�L�)��}TD��K�0��%��!�|����MR|�d2�u%��Z���#V����
���Sh����'��t�-�6c�0��B*{	K,;�����k�8BMQ֖����4p��� ��H�'���Bab=-Y=L#�bsN����[D�Z�>��P �`b+��󚈣o��=��d����r���֘{�ۆ�Cc\��[Ms	֯�E���.G�?v�u�y�$v��-I�z7V��/�]����h"�"��7�p,�)�R�^t?�3���U�\Kd5o1;���G�����ωGb%�e��Y���Kf���^��m���,���)����T~/@�ĳ�^�|֤g�x�rO�|���4�	��jq���w�卹��%l�l,a���*�>�`s���JN�>P��T��F:�F9���kǊ̳q�B�x�h�f{��.{ܾ���rð��Bc�4ܱV�5�:Ӕ�A��Pc� ��/��`{��IW����rډ�2�P�y�ǉ�ri0;��1 t<,�C�P��/N�l�J۟o�T��q���)y��$*����=��c������$�4I%9�Cav2�� L���պ�/Q�>�3,��R�m�5̓��&E]�΁����Y롢>�����l߰�D�����D�P��:E@%(�ʳϻ,�F/�=� �GrP4��[zCv�K�\�4�RE��B8��B}�N�L��+;��շ�zG��̛�_)��]2
������켑q�E؃G�|�c�pk���_��,MY��|�]���B��F�*�����8*m�~���EA�	|���:J��@sþ 2T-���L�r{љf�%�8�h`IrAރ�TI`�"̚�ћT��p�'�T��##�_� '�A�"�����Ϫ�w� ^@/#l(	x���$�kcyLiLp�}�*�Z������):����H*�����q}��M�4�ʤ�oZ�ڒ00����ơ]�!���K�b��B_Q`i�+Qp�Jq�[���mb�<��|�F��AkFS�@�����S#�����jM����hO ,�?H��8E ��p]�(�k���.��Jl��_
��E%@f 1%�M�O#��T�d1�d��Zp��o4d��q���a���g�h�q�?�	�y{mɫͱ�����'�
7��#��بc[��[-�D����Z.S� �]�u���ԥ�d��<��hk���zs�X�:���s�H��m�����z��_�M���M�~}8���?(sk;�8�4�;%*N��E�rT����0�Z�$�>QU(�[��=�ܖ���g���}s���qI�^���JkyH��M�^2G�ȸ���0@�s�<Ґ�����BIBQ�>e�x�\�4fmd����BS��aX���t��e�N�w��W�oľA-��9��.�wX$���a�@}�S�0���d�o���.�����~�f'B?m���hƍeaqI^3�a�N�v��鑎�(`��a��� 4CH�J$���u����7Ɇd+D/S�]�3���"D�����F}~��h�-��t�޺˱�q�jQ�z��H`j��
Z7M��Y�����)"�:	%�&y9�b�dy�WF�-���1��}c�Dw8�&���3�gc�� ����63�h��O�y&�u�����}a?�96��۪�S�ݑ�/��Ei�[�����B���tN����k�<�ѕ�ٽY��0V��D<,�dد�
�5�i��#4�P���r8�>����ɩv��FP�zw�ω�P"�ȋ͠1Ӵ,Pņ��(CO\@IN9	t��k�ĵR�b[wy�z��/�CW+"�9/���Fuq��PS���b�)/�M�7�O(hw  6�4E��n2���-Ž�/7/�NB(9�h�?��=*ldn��L29����@�l�_2!��뇟�CI�L<���ާ�"e¹H��ys�<5 ����V�q�3����\��EѤX�ni�Xc�2�S	�Ohm�1N`X���hR��z*�qP~�x`�C����ǿ�Nj �>�YēK�Ro�4�,�����R����$B�"�c�;6��0��J��u0~�}�Z�{c$��G����*âj����Hw�<4HwK#R� �C���!��-������������w���Z�v@�ގ<�Z�ba;\��2�JK�p��� Gn/����� �F{���[mi�ZE,��8@�����~�"����\���@�Xb�����6���� �3���}�I���c9��h�/��� j�B�C�J:�﶐��2s����D�Q����]4CW ��xc�|f��Y�1��CI�܂���=�i��ω�,��h��nn�LԷ�B�t�����Ĩ?K�6�e+4�~H�1��� ep3�RO'���C!](�(Qt(y����,�D��JJ:����<��}L�
g)��F���N}�����y�c\�ss��c�L�J*s�P?dr�[�D,Y�T<̫���Y*�>C��Y2��ŝ�_�aW�%�:���ۋ%�|�h�.[�Ǟ�L�"yx}�l+�td�	Ry����aVх�?C^ P�Bo�_g�ҙz)����JM*E�r�ܗ��RQ�o��՚	�ȃ%�"����q�h�ѳ�4��0�,P�:�L�Ժ�����ko�
ī8�Q�����~g���L���b�>��@lқf�pj�s����/������s'X�LP'���яƝ� ��_B^[ݝ:JuD�ؒ�pK�@�Uk��P���4���F����$�oK��{E]'��T%yM�cy��h{}B[Cx�F4p���`�yE���8!�ó��ʹ)e��vZ��p�͠�r�Y�8���	��)Jr�G= �@H)�Z��=Z� �:PޖTR�@t6�:�?J-���/���0�������Ibi��E_8uMBl��
>!��3��2��I����f8�\���lB��6�#��g�R�0���S
�'7��ru�r�3l݆8����G�9��f���n�T�gJ�e�7�鲁�����+�TmC�8�q��Z�^�b(��-|����Q��X��tתJA�g��ܜ*��) Z\l:g\����M�tT���VZ@p~�u驺��%ʡ��4d���kC���m���%Cı��Hw/��*8nG�}���i�P�Z��
���&�&�>*�ryDLU#��p��[�@^�%�����O��\.Bj�VMM�-6����r���yj��~oj�E�1��S�$X�m��b$F:v�W���rw��x���Ls��՛�t����%�ƥ�z�#S�6���p�6C���ɒ`Id���jg�ivQ'uuZ��������XCc'�X�����-���:..Y����r�󑗴�<�2 �=v򝠳�N��~畯_���	$��sD�i��=q5rJ*<�K�vw˥QR�)8iq6{��VA�Y"u�/f��R��~kZ{s)l�e��V�
���FP��K(U�C��7�C
����D�GK�b��a�8g�B����:P���|�v��%�U丨��叾�,�n��%���1�6ˁbbY. Y�UT�����ڱy�ꚗ�j�,C7��hE*2�K�p/�d��:�^C�;�P�s\HA��npH̝_�j��t����y���B$Z�0��7��,�[<#�x{Ԝ"�����w���S2E0v�gpvʒp��|��j�M-7�ҍa�F7pu��-'w�򳬌a���a�,\�?Ka`�f�Q��r9.��#G��(���m`��T|!�˺��q\3k�w�6�>u���c:�s�͜���9xB���p��v�G����	ʦ�:�qv6}m�����y�Q�f����M;���41����%5�k�z���8�Bs�b�Id�����r�
vĭD�;�~����I��Ze�R<�_N��]i�T*A���l'�[�F���^�Z��Lы�ۿ@s,�B�$��;���	�lkv]����Oo���9�5�+�/w�S�}�M��C�e4"��
�FlKz����=a�2޲k�v{�stq������k�<�m(c�~,M�i�ٯ���1@�d�y��Z1AAU� �V?WrH8���Ԣ~������1����U_�Oϙܗ��lηN�?�zW�x`Ɍ+޽8x��<���U��Ɖ'hk���W'�s75ظ����䁯��ݘ|øa�� ��;���t(�84x}�-��cd&�8B�n����Ku{�(�&�9-"���Jz:��Gl��<$4���'0����7"�c'��K>S����˫I��%K�{�`x<Q~c~׽)���B��wmΙC��/�#n�[�<�i|��=�$�y���X�PI�v������"M��`��``�*�����Lm����` 1���]z�cҽ<d���[��@�j�����x5����g<J�G��ȥ��~�E2��ڼb�'r�LY�OE�:Y[���S��_�[�m2���h�M��چ�卣ډ$�� )8�v�Qo���t�|n	2[�`�ۧd�*Kk3�+>��΋��ǳ"a���,���ѥ�.��-��#��.�1H�	m<��g+FcÇv����lwjq��\�.�̜�u"�{�J&B2^���K�u"w�Z����R����]��x�G��������	�c�o�i�e�I]	�wѸ�!~D�46kw�&�yr�z_>�.�mEU���+�����?�䄎�/��]�(�o汦�<�C�)ח�?D�܌��a9��Nk��MU�P�.d35�1����j�bn\J�Ĉ�#h� l*L� j箫��X����]��Դ��4y�J���9!R��Wr�����*���keȹ{�J���o;{C�����Sq��Kl��z�Q�sIf��ͦ!��"X>���s���7{�i�m��XIOb�/E/���Ȥ���g��i��ɥ@���t 	;������h`���x!����]�S���v�C�u#��"�_i�M�}<z�_r��$l���L�_V�f��$`�OǾ#I�q6-�>��9�5��H���Ŀ8�K����yyGћ���`������|zg�i�~�����*���S�+�!��v��F|x��Ŧ]d�O0o����/�Z�9�QFK�W���*��5WU.zwr�:���ad
}q��.m�B��G~��@����l�]�'���r��;x��@��u�:	�/�B���	����������G񣰚5^L��+ݬ�s��m�`��D�4�L���0k�aB�;sQ5�1&�Eʜ]?����z�����:Hb��˫��^S��sB���2��>理��h�����0�8Y."�-o�,��>��������2�����-vxo˜��#L���3Q"[A�^s��0[�ݑsH�Pޫ_�q��S��ynNo�X�n�/Ǐ���M��U��N���D���,��Y����;p�Gmn{��K�F^=���U��X,͖qnU�m8:d8�7��A�7S��乒ޓd�pV��	0���2~�]�p��S;���Aa^>��cZ`":$�?d�'�c���Z#�-�ܰ����0ʑ!���^~ ��bŤ������������[3���MΥ��S�[�����*�j��xcG�%�#8*t��@Rā���07�����m�$Y�Os��4�V��W���ҜEw��L�aR�PW�#{�0�g,��ZI>�Q���Z�Ne���X���~O�(�ҍ�g�7�Q�H�g� ��Vҏ5`����ǥ�)C:�ۿ|k�� ��m����4�+zܧd *�Gl?r{]�[��Q���^�ҏ8���m\�} �l���tv8��+�扙.�@Y�u(j�-;>����O?u���9�|�a�Jm�0��0F�(��
�2e��Zƹ���?<�N��I���ugr�Euv�e7����Y�&��2�~V̾`UN��-�����
Ga���e�l~S��k]�S�K�����>/>]Җ	�}6߬�4dsϨ��6L�Ǿ�>���r��U�~ɯk2��>B�vA����-5��W_���,���u�zT��k�����6��	��� ��ʌ��'.$c�y/?F0�v|�=���i���q°ed0Ե|����-�0�Lp~�[�~\��`�=�hQ��{[��ȗ�~8�����!S���]���*9ӌ4�$�B�èV5��O��H����:�M�A�zB�����������+�wANry ����4��wr��4E��76�*x��PD���F ��j-�?������E�@~n�MXWA��g+��
��J�{���o��&xA����~U��+!&�~R��xɊ�Y!�\JNʭw�M&}}=emì�<djy�N-M��Ƥ��y�
��jȍ�'���ɮ׫ڑ��(�Bsy�H��qU���<~k7�|���ģ�����\0�|m%�U?{������l9s}]"м��%E�b!�:W�/5���͜Ρa׎���G�6�A���z�ơN,�������"����="�7��=�+���U���(�X�Q��*M��w���ֹ	[Г]�^ �V��0��5:������ �v��W���XI�)�T�����"y^Ya�a��³����Ǽ-q�ߖ=8����P4�����2<��H4�L�G���܈�w��~)[�k��A ��fw)���Ǚ����;	��O�@p���}&���S�o^Ա?,���gyx�i9��mr�M�����cP��$��$k�����R{� ]��
d�]|y�k�y]��*J����ʱo;b�[t<YPur���jVR��x��o%t��*��u�����(uIZ�9O�,��"Y͙�E
2����b��e[>���^(�щ�2��)֍h��_=�V%����hv�0{�������Sb��^�#�,��b�k�TϷ(ȟ��Y>���Ց�F�����1�l��
=��;o'��<�]�9���QV�?fC��[�#�R�������2���Һ�?�-����;���A�ɽn}
���>j*����6�O�OVX6O=��{wf8�P��=H=���� ��K^�9!��T2�~�f�N�u�2T,��u��r�!�u��e�a�Ur�'F��;�B���/3E"��``o6~�w�8���~���b�>8-���(;�_Z��H�:S\8�!U����Ȁ��*ۓ�@'ʕ���f�Ҙ�&K��G*?w�J�дC(V��-����1b�FCQ�%h�tSQj(�
��o��_��6�y�_�Y"7eZt�jkձ��++ܮ���b|�&j=,j�2s�^����C���<dG�㦕�HX����1��ڔ�K���'n٣Z7\y ���������Q�J�Kl�@c�-�'�íw�>�=��Y�%�W��2�l��YD_0#�W��/_F���+�
1#�_?�{�=jaӽ\���"Q�$���H�dW�?��n;bX����	O=�u:�^�U޷v��$�B+ʲ���=�����������ƼP���Z/�ʋ�U�N��ELR8�fܟ���x�ڟ��\z�u�?0e��YS8p�]��N�]��`M�W��
�h#a�@%m��^���L����}fz���R��O��e�c�4�x�$G�㙲��N�9T�b��B�,�,�x���4P�7��6��f��:�v~j�F廘�"�ҝ���ƛ��c�n�Z`WAJXe�l��a��h�����fb�����-��3��U`��?\�L���<��F褥���!��޽$�NEC��!鳹�2�E�����׃�',�L"L8�K�xV��x��T@��Q���K~*��J`7~�r�!�����|�B�r�j��5o�k���Y�/.�S�Q_������D���M���r��,k���Qg�jq���8N��-6j�	�B?�Λ	���T]\�"��
�R���o%;�j�o����/�W/V&2]�g9Ռ��[y�^�4U?��>E<>�Wk��&ã�	�F_��d���f��!�l� ��SA �@J�3sǉM���k0$�����Z[0W��}��O�A��Θ�v��Z��SϗG�q.�GI�g�j&��:�P�KH�P�דcRO��+�����1i����ܻoP��!�&�j�j��Dx��Xv������w�!������U=m��VtkZ��C �s�ͨ_���U?���VA��[^�d�._5�ˬ�D`XW��Gٚ!���r�+|��B 3��ͼnN �V���,ʟ.ߺiO�EV��J�d�0���v5Pg����(���=��ߐ�%�{�sz���d�K��r?/����}Sw9�N�}��$�e���>����g��s��Z ��-6 ����ѡ�nk??�?A��Uk�$ r�yQe$-\�RM�M}3WKYH���_Y�X�Ω�E�6h�Td��F�s9�W���?��7n�O�aTǥ��#q��]�%b��-�K)'�<"��"��=Ef�P�����_G��ʒ�h�j��
!M�����#�s^��M��X�ć��v����E�eb�ҁU+ʃ����-;	��́�����>�}��6�U8��鐰fߚ����S�?w�@Qe�}�x�l�罢��p>(k%ƅ��L^_jЫ��.C�-O(?�v�C�,�s��uG��Yms�o"s;N3���	��^�8��9Ujm{L�/�}�SL��g���������@8�C�y��x��<z��P��[ȼz�lO�qt�\�����L�ДZ�������2�LR�<�L���mb,������cȋ7�6����%���9m��U���a��)�@2��e�G:�g= ��KF,�+�!uxc�����z
D�F��w��;�~�$��V�r}�@�'��}�����a�%��Licޑ���^$@M���2�ϡ�ˏd
	�y�=��U��u���AQ��p�4��6�p��9d�'��S���_h��o��X96վVd �4�@)z'Q�D�6)����"�%�[z$�eճ�z�7����^ܟڜ�y��i6�JV��<k��7T=�]0Fr�����#H+C�k���
��R� �$�ݘ�]I�Y�K<��(?�s�S��3�gp�Ƽ����",rw�S�Z(�����u�zP)��k���Ĭ�6׺o.(xe&��=οQ�ss˝~���n,D�4>�:p�	�a�~��W?����l��Rۄ�:�Š|9�+���dSy��X�����
���΍�>��W�$PVt�_���6�I���Z�pz���ؤ� ��E��-,�?��&b�u��Z���^
�*����̈́��9l�8����O�o%0"	��k�by��hck�q�4�C��<Nvt�!��(�$<�F�ɰ�#�����U:>����m\�,q���P�46	�h#�&<a��F*i�ʌ�$�"�4���k-���qj�=a@�GU.33��H-?�F�9�Z�O�h��k�+^\�]y�lɨ�£(M��Ǩsd~�ͺ%O\w���D�������1�`5+�F�����Q.F��7"��a�d��yj��KI�!��$���ԏ6������|'W_x��/�($1nt�X���1BY`#Y�h�O��(�W?FB毯�""�:�J�[������N���z>�ʵc
���5��i�j�1�+o�iPb��=�OY<���'�CRǏ?X�����xq�=���-Ѱ�1n�Q�}���/6|VVM��i
]ֺtc�[�� S }�%/o?�C��d�{��Y���G0���e��g"
D�SQ�����agݐ�R����Q*I�ތ�X��^Q^"�*9���}��G�����f�Y��XP�,�hty���-$଎�Z[���,�H(JR����G���&�u��gxo�N|��
��5�ܕ��b�2su!14���_65\���"6�87��a�<o�"� ��u_f��4M����݀�,A���Q��U���(%b̓Q��_W�b��\�0R�������ne����c������x"�� �M�a�n
��Eok��PN��O�����m�b3u!˄�GZV����D9#!��'���Z�X8\H�HK~����������v�Ӓʐ�����":\�臤�=�HO�q%���ߵ�2Ʊ8�#��Tz꺿U+�)I��a'M�{��(��?MW�R��2��=Ɍ�#��P]|P~\��Y�U_s����p?����&�-��֡9�`���:��Y)�� |�G8�w(Qw��n�:k{�a4;���)朞w��j�(%di+�m/�`���oi��lo{�lyUr���tS�k�W�Պ��'7'�anЧ�m"(�F$\L�,��vj��X�W��k{�LU�,ɨ��Ct�����[��Ĝ�q�kZ[���.����*��m��O�©��%���e)���@�X�i��`@3T��h_�����'$��ZB�ّ��o����?�x����0�%z��v)A�pA�Z`��0��i��VY�1_�0z[��%X��x5��\�3��o5*�wx��Ƚ���	a\��c�qs�2�������Nĩ�a�gN5ߎ2�4�G�zo�������V��6{x^�Ώ�F���~^¨d��������>������VݶbN�s�&�����G,_�K���מ+�����L�ٓUP����F�@�3_��\�sW�R�c/��CV*�L"Eޘ��>��g�1Mc�q��x�V���!T�n˜�liO.���*���yWiR��U!���^�+n[�u��Q�2+	�ū�k1�Z������ؽ@{2�V>f�Y�>���f����#���X����ͨ�-Z�1�Uw���[H��X1�����޹��n��n@��C��4�z-9@����Y��͑�f��N3Ld�dn�R��c�cD8%���#�>��:��ia�W��I���[�Y�6
l�j�Rn��)q������JrPq�,�������}ڐ�F]�c�P�XOS�<�s�3&���l�5길@��OL�5�^�6�������k�R^�xFO$&'�a58v��k����He�2��)�u?�=&�/h �\�f�H� ���Ì�$��Ȟ�u���������M!�6�Z�bT4�@q�BU0��]��]e������2��������ʩj
�&�&0����+w� ����R�C����wN��!�7F/)3'��3'��A7l�h�'fM� :4˨\�����~l)�����rԧq�CRZ �I��ȼ�;p`i��-�4	4����Fvٔ촕�6��J�#��Z�`[b��ڶ���#��H��K�6J�I��:�����=�E(�|������¯�r!�-��+���R��8�~�\"�D�a��p���%f���H�u��_:l�*�Z_��䍲���~XJ�C��q׃���b���~�����IW��� �¨0�qDb��⽻����D�@���%��+���h[Mz��>��t�����xL���bS��NF��7�����y6�#b�e�`�̶�u����y�( ��"��'�ibz^�����Qz�eFcu9pX���T��*�̾��e/�~\%��������
�
�VJ�]Y��%�)R|���h�*Y���c,|0=�����{	�CB�r��|��$�G* �n���o\����$f,�����뇆<.#��F��YY��L�,��f�\������Rԋ�ҧ"��j�)i�Akհ��a6R ��D���oKL �Ɗ�f'�ϫ��A��N`STy�v������
?���_�p�h�AD�|9�<�����Rgc�0�ls\l��U���m���  4���O�Ǘ�!�;Mr`@V_V[U�v�$�?��ɠ�tp�2�e���k�z�<l��9Ϧ��ܴA��td�Y��	D&���@�4�"K���XS�2������M���H���9�|����ѭ�;�?����LJ&�CMrY���3�'����y�~�p�����%h��K4W��O��R��;�z�v�e�����`�Sql	�<Ӳ�ߟ8(�̭8=zHyJ�-��\���*U��ɖ�z�څ�.�d������y�����,P�n��c��WR�f4~�u2(�̭��9P]��� ���-t�m�w�MU?�r4��$����v����.�V����WG�K����{`XbZ(��p�C�@g���\!?�+ΗF޻($�~�^#�Bt�o�vr��M����JNEF�Rc�*�?�;����"}j[���c�hh���H#��Y.�>���	�ˬ`��t��ț����d�����"ϓm|�J���R%�ue����V�|j'�t[_�dY����� l�旚*RvQ���P���� U9\ݨD�{v�K�6Kďc���5� �^�������@�D�$���/���w2�����G�g ��Ȯ'2�����g�@� ��*�6�Tn���^�뚣g(�������DX���v�eH�wQ(E����V� b�n��\Ć^м���gƫ�Q��r�ޞD�ݕ��XT���RXѼ"�����Fa��ߢ�M$��yۙ�ի�FE��ew|���a1:\��&L�k�>�ѥo;�(Iy�M4��6T� ��]1���>��YI��
�垈�z~@$Z��W��I��]���iy?�e6�?�h�"�큒��p���?G�v	a�4��XF{�+��9�Hf�sŔ���ǂ#*���;;f&'[�v)ʐ-�ƪM=�zn=�yV��i@V�20F��9xt�PJ��Df��Q� 	{�.����*��S4>�Q��ޝ�h�3;�>d�5]�O�����}��K(4���Eyt�5T���4�����۴)���8:�W�-ޓ��v;������_��d�z�z�&!,#9�&]���iA��T��aw��U�������YJ���F��+S��X!�Q��3��߶X��b�u�����AKq�5�o=��F���B��ч����[��=U��?��E�@i8jm[�,"���*R�O��H=�!Omw����U�_�:'���b,�L���	�\��\b.��Z�ZU�M&�=҄6�7��b����q�Z!XږƵ}Ҟ�N'
 	��oLn�@���� �tΟ��l������c=I�|{M�j)^sӀ�	�:����w-bK@BQ�E����-�m]�5��͕<9r� l�N>=���1�݉��C]Q0D�ř]Q�����+GvU�������Ú� ��8Y�K����G��׍w�<g���2����_�
�_�)��`�׮�n�o}\��@��IR�`M�����+�[Ű.^���Q����x.,��C)aQ��K�K$��������{�(����Q@�>���|�_����@�3�t��V���n�jJ}��٬�����n!yӻ�u=��Zp��3I����U��*��?U�e��S�1 �R����sFny���������倓�Lv
b�&���+���i�G�~��G�zα��vҠ]t����$W�g�_<$�*� ۭn��k�=
����v	�D8�7��b]�M��In�D}�.��C������L&�N�U�d���&}���,-5l��C�Z��'�	\ �@�[zAihmDpC.A�Jؼ�m������R��`���e?�/E}9x[2�:J�Q�h���rT6��D�������~d4���u'j��-a�� �O F�3��7��_ݑ��U�q)F�����uE.�ah��F���{�
��W�4�$lk��$C�F�ev_Xc��~D-E����YHK�|e���Gü$�B9q�W�{[���[��*��НW�w�Sz1�
�۔'�P"�R�Zt��������6k4�c����:�`�ϲ�l�@��('����tZ�~��0�ʻ�BX��s��]��Ti���22^�w�VRy?���"��&Y�;3��Y��Ʈ
L�{���}�6��2����@͇�۱���HB�_Jv>ǃ^�b-t~?ƨ�GP��Q����5�M`RM���**������Y��Tr�K?����	��a�#�V�΄�ͫ�L�~����U �T����ߙ�E�1T���,zw��yv�K�.�����P��ÝC���K��`��s�s�;�'�G�Il)	�����o���&����8U���L��/L�H� '	d���H�I�1���\Jz���C�T<��;�������K8�bU�8 ��7z�#0�B�F��M�xDq��>l9����s^_~��:����͗$ȇ߿)��q�P�V�y�t@�T��&k�?�T����c����������x��oP��i��6�$�^���D���bX���?Ioc2"�Z��/Y��&%7t0:���q�PY�wf���^���헃(QG������o�H6s糖=�^��\rpF�5�P�w�����q9nXe`��pY�r�P��y���4���ʀ>5iz`��"U��h�5��QI�!](�{�_��Ð�Д��׿�P��
���YmNx1�R�lxxG݅_e;e�x���ًT��J���@�d�F�::H���h��L�V�XL�0�ęd��]��I�P��[8Ocs���r\L�d^H�o(�ޛzT���X��5���`!��RS�<�#��I'^_�+�T4Q
��v{H~�����O��(�u8��qL��,7�z_�6�����lx8��,o�z,G!�Pr���]�bF��s����DRө�|ù�c	��|@)�Zw󾽖�&�S�U{a�q{V#)Z������HA��/��oO���qB_9�u%w�%9��x�ft�5}����f�۪����&ƜoZ�P �d��Fv}�O�#?��&6!q�$$]@eN��;/���QG��JP���N��gj��6τ��6@EN��»� �����g���-���4N��_

�L ��o���7s����	*O�`��s ���x<�>:�"�����1�se�`S���ݤ��l���G1Х]�)SF���~z��H���n�ïh�$�hO}@y���>.i�V���M�Z�h&+�</gF�dJkЛaR�l����	3�pI�2>r�~�z��!��2	�+_�f�^d,̞qG�[X��}�nQ|J�6����b,ܞAOtsx0�/y��,E�����GH9�����.������ʘQ���G���7x�-�j�Y�U`(L��3�v�<�xK��,
M�	���a0/��-Z_����w�Y�&m5��(���4�9�Rv��g�o�ovL`��������cz���x��r{�̀$��7��~�L1�V�S�����o ��%���B���,����	A�Е�N��6�?�������ǭ���r��i{���P�Qy�Μ$l�	�����Wbc~7��k@X���)H�N��LM�'R�F�Lp\�� ����<W6Q��p�l?Ѝ�`����'�@=A�j 3�!�4���z"s�D9AB���%9)٠-�fܿ�jg����3pSG���U�i��F3����JoUU���=J���F����/aX�;gW�BiVq]^ѵ�_[��m���P���il�N����$6^<Ѐ�ⷧ��>��jh�$ �
�>���˙&rYQL�~�Sk������!O�R�_�/��� ����f+G�Z��p�sW� ��lސa�v'2�>5`X"4
"3���H{/u��j��& _����Is։�@R����٢�J�a[i� �(��^��� �����g����w�5�'�g
�F��R�p��K	���N!��`�'�y�7�yAt3�?�~z�*�����,����o��9�+n�O��i݊�P�1��c��К�7,iԬX����%�!@�}�lZ�\J�����~��|V�q�މK��䝷�"�[���.X�Z6F.��a��?����q��&�(��҈8���')r膤�|���_�Q~KX��N�$.}2Y1:V��Մ�uO��0 *,�H��/��
�w,j��P�lIYcT|E"6�U������`�03!b���jI��^��L�ށ�$���#���-È���ɟO�ޑ�&��{�CK/v�,a����~w\�,�
߶���o7�e���ӓ0.�Q�bu��,�%Z���y%��2n�~ZBB*�� *{,&�����86II(D��k��e.$��g0I�`rZ�cQ�H0���Ad��5_8����P�k�Ԃ'������!ڋbЏ6!	~�ڽY��u��<�)D��R�fU[&'	9+"(���G��q"+G� �c�9F3�F�@8��4�����s&u����@h�L��{�|�}���e�]V�U�+7��<��2#ʔ��U@fh���ud�W��6hIe��{���Q�ŧ[A�逻��(֌�����<$�Qf��GЖ����[��b:��*�0�p�����w��#���.�W�b�1�a("�M�W5��E:�.v��`%�$���I�5����[`*Q��l �q�ڍ�:�v�T����p�ڣ���p^�0U��2Q?5B��-��n� �|rB��g�$#����{�?)�>?�$��� !OBW��a4�yR�yV��B��u���"*��-W6�ݞ�Dz��v��7v�#4��y�1 �fm�o{������_�1��E*^[�o�r�ѽ������S@��F��v���3��8o`<���Q���W��؜<Dh~���U��������<��{y���)��sGD�S��T51۪5u�D���Ƴ�>r����Q���F���(&�lF����'�+�Y����E���`��u�.�֚���D��b��x\^���+�{��%s�/�<��Eid_��;R7L�	sR&~�^l6ڨ	,��X��ۛ��WR�p֔����U�A��oI��IU�޾�U�%��	�fw�q�j�+���p�[���Kº֚-
�"*�6���me��蛙�*�I
D�S�/�_ ���,�!����7���XD��G,��>����� `��gW�4	t���x��Ǎ����@H����!�Ϡ�Y� 3�_�@Lp�gw��GR2PM"��R烬E��
���b� �ɽg�9m2u�<�%�q�� ��F��? c҅D�ꙶ��$v�����8 �i��$���b	�\)"�C�Z�X���Bs�]<m��2�I�%�k"��/.��� �f{���z�1i���.Sp.}��
�mD��<��) ����Pf��X]��i�`
�� ���^�P��~�����ML��n�����K[�(W��R:��YƚnÛ�e �V8ߎ�i�4�͢�Sh^��T��_!*Gi7�i�Ξ"B����}�r��K����/���K�*������Q�K��o3��3���<av�_\qq��w
��O�@�风ә��a���Md ���[q�&����ʹ���Q/Ox�Kls��gr䲾��L����j-�q��C��9�����ᄺ����m���;�(Z=�4��iH�ג61@�?��| �
q3S�u���}[?����.��x1t?v�gj�V���n��ɒ|?��a�ط�m�4c�TEvr蜋G9�ng�<A�^��Z@�qS��^��T�)��w-XSzd�,?z¹\��i(,I-[�ȣ��@g��ﾲ$���06��#��Qlx���:��/믫�F�ާ����8b{�a���,_��u�il�����n6]8Y�t��E�Ѹ�Q����IVD�'*g��8�(%�(7�N!2M/�R��C��R�+����i�z�����oˊ˝Jf�����p̽И�c-C�S3�
����2��ܫ�E�Q'x#�>�D��g�j�{��%m$jn�kA0Z�vjE?1�+քD|^��y]/����"l�\��R�.k۪ASO��Y�\ݢ߶���+�i��D�Q��Ng3�=<�Ls,�ڶ}BQ8��aa����؇��sF;���dr,v�?��;ޤ��(��wv�+��c��俟A�&�>���C�ʲ�k�M�D�[���Y3n|��=\���H4y1�&��k����ʢ���5��糶�'v21Z��d"9����}M�Q���򻒪��&.�������n�5��KyA�@�.��O���]�@����Qm<�!�-Ĥ�̧	����h�eCTb��Gc�T=���k3 �_n=%�J~���z�5�}$*r�؅A�=L�����K����IJ�ٖ����:�2+�x:�썹��c���o�.I�|z�W�R��p��"�<���4_hR:���W�,!��P�m���*����w\�=�6ٹ���"����P+bW��LJB[F�8[:����T7OK�]shv҆� ���[�mw<��g��4��6�f�Yn?I�4��e2(��(DE�QU���H%M�v��b�w.s��q�h���DN�u_@,��i�r�JNk�(�g��y��J:$z^��ZL��r�`r�T⿉�匂19*ۙ�c�ʗ����^n�V���i�j杰�n�ԫ��fݲɣ� ��!�Nkƙe1Ӿ4���W��u=(�x*Ų˲�I)A�h4����n����@Hk3�{i�=�p��������]�|ͤϵ�a�/�Bq�\�]5jja&�o5�l�=���gn#�Z�&�Dj ��gmRD�����Nę�����#���j �+(ИY��ʮ@@:u6I�9�RDn:���Q����w���1�X0�"V��ļ���̈O�����=��!�4a��<Fbi��z$�a�7	�-/c�*��	+g��q#���/� +sV1����ssyc�l ;���S�C! A������Ig/���R ��1&?#h{��.�.- �<����{\r��+��%���i���c[�F�	<�`���'��KN��Bpww��w��y����f�ݧϩS��j�sc��h�CP���2g�����7"]�8]%o���Sj_6�&H�%�P�_`y�k�=�@='O����Z*Z�� Ś�g2P�{�5v.$~a���2�^�m�f�������g��Y����F �U�K3_���������$|]�-�Tj���
WM�kd�|����";�o/�H�~9������f���o���L�6L�H;yj_��\�-q�k�j<����`����m�`�<���3������;���rY�M�Pn�6a[9XFE�ޙo�]�u�o)�] �Aq���{�+�� v(�ܜ���%���}��!oc���������WZ'�z|���zC֖�Ҝ�"�zϛ����·:��A�tjmev��Ӫ�����_`�)����� ���F�^_->��Es�G���~���$��˖�)2!�F��;�dZ��9�̭QY0���<����T�<���׵��D�ї�;��rх�HGv( �I���a	�YY�2��+�K��x�驋�����I�JӜ�^"[�?��w޿�cN�Y�upH4� �/(q�V�����`�hqPd�캫�=ws�~2�>-�}�����rQ��S�LL���Q��*ۇ�U�vd���㶋�p�U0sJ�*�,�����F��f(�a�]5�6��7�J���#��W�w�H=:m#��ߊ�h-�-J�JW��,��H�-�̲4o�F)	J�j(Ye��zj�����!��s،E���f�H]�T�o",�Tf5�ƞ8C���D|����s��Iy�w��q�:#� ,��o�Pw�^���ퟗ�����j>�t�t�v�[y�E��8N_��ܿ*� �% n]����ڬ:��eD�m&�UG۫�LB�{�:؎����$���Q�zw%&T�m����K�~�
�x�q6���ׯ����+��� u�xLĹJ�*O��4{lU]Nd�aF��!\�7"�T��6M{o��à�m;��c�1%~ke��x-
�b��K����������F3V"x~�i�x�:�	���mp�$6б����P�	ެ�z��C�X�cZ}���*�d���n�.g~�K0����,�I^�8����=���3h
zt�.�jn��n��֦3�jtMAf��u�e��b�H9�V��7Ȅ�*e��'������̑�=��l�n�*>�L�>�L�d�<V����~ɥ�Xl�w�� �(�Π=���FY���ӥ|yo�b��里k3Y
�زq�_��7{~��8�f�\�;�ǻ�]��C���|L�YK��贉k<ɪ��I�, ���~�M��s~�~�4��ϋ�TetY���Y���6:C�ݶ�����?�?kx�0��h/�*n8��Kw1�E��m���g��˪A��g�/|���m��C���H0��!t)�qp�VEm��Kd�v�a�싟�	��&��
��J:�zz���5SH�ns���>����V_�C<7�����;�Ef掠�H��u�)�ej���,6��v	��k_^����r b{�u��/��9�%쿛��M��5Vm�h��"i��x��(�:C�i��.ج]+��%?|��V\�]@��~�a�f�3�w�Z��ۃS��'�BǙ��gi�l�������j�"�Q[�Ȝ4��\/f3�����q�-�	Y @4>��&�0�{�>_���{����h,���y��m7��������7vh��U�R��J�����ui� ����Ͼ���9}$7v�@3�J��oZ3WϢNe��خm��}8e�ei��g/��FDq���彔���/M}D�@L �}&��������_��BQ����SJ06�FU�ǌ�2��J����'j���o>�e�7�Һ��6��Ԅ'��ɯ�Z�疋*}6��g+С��x~�u���.�j	��/��i�s�opH�o����?OưEkJW/����I\�u�S��[��t/�U�<DW��tls���^����߿.��)e�2�I{q���{#H�:�1R
r�GA�%��Z5E��}z[���lj������]���JN����ifϣCH��͓ݾ`�d�w�kt�6��<�#��e�HAUCd^��I�*	�,�'�E�]�/+�7�ή�ë2U0ɕ*�����&$"���e�%���f\ݦ����Url&��'?xM�/4^m�\9� uA��p���#����Ύ��'���2����W�˃��>�D`�ZF1.g5��ӽSz�Oq53�l�%�c��C�:,���@PevL����(��PDjPI�e�cH{� ��9��L��l�d8��������r�MUm1��Q.�z���q�?La���+������m����dPk��Ul������d��k%�ZJ{��������Z��6����D��O\�1F�[�G�}���y�ƽk��8��%��Ɍ�#<t�N�����k�z��_F��^Ʌ�*�o�A�w�-	=޿��&z��R\��"Ɵ�v�\RQ�ϛhQ�GS'`�QmG��T��������������)�#I�`�=$���I�;����x ��d��!���,�ӛm}u!k�T|�|�;z����f0f�޽Ǟ�s���&2�UZ�G�R��8����-��
'7�}>3uVG��Ċ��z7Z���
�Φ_��$D�Zr��4H"a3�g؊�8��z�G|di8�+f�L�AH��<�ag����]k��Q�OX�aG:j�p�:D���iQi?������e_�a���VB�a�ΐ]��;<9��7H��9~Qn��y��G����,�`�文�����r��:)��ר�a;��۴��9��jq�L����n��v6j���g����O��L��i����|�i�{³��膲�}�j�F`ϛ~�q�M����<����܀�l;��E��!��yCz����JD�|���G(C6Kc%���gΟ��׺��܋�����N���+�O늞7ɪ��[$!����%��>5���q�;�9E�G�o-&���m�"��"K��_o���x��d~��������� .d�l��Iծv��X��R���������2a�X���1�"��T��d�	!yr�j�ɷsN�rj�e�]�LH����v��h��Z�_7�7Tt�g��I�4:82�k���(T)[T�)˴nv�����������<U�?C�g�K�[�~@7
l'���N�6��t�NciG�F�g����R�B�f-�%-�\��+�d�m�.��$��@�5�Ě[)�X��v>����h]��=���- fB�5}�;	�<ͶcDO�+Wv-��:.e�R��`M3�l�j�OxF*#������V���\EiZW��屄_-˻�T�H��]2�ա�_�����_{��@���
�J������X�e�x���D3{AU��daI}?Wň�������*�f溒�G��}J�����|n�Ͳ�<G��)���U�Ōʖi`TEq�3������������pg� w⟿c��G��&Ï�/�A�*3�j����j�[;)��1��
>�4����ǨO�Z!�a������t��-RS�7�l
K"��@�?�I�.B�}�d<�������������&�r�a#ʊ�B�ޘf�y�c�W�BZ��aweu�-�#�4�Ś�4�~>�8��H�dg���q��O������U��>��ʶ��W�����63�^��t�C��v�~���u�b�uG��e+=<��<����V�n���dlZ���y�%7|��8�`�V#�M���"����߬�$�[�P�mz�Qy�8��_��BM��ww��������,����vS7�R�=�XcG&N�E��4=YqT6 �ɺ�p�ヱf�Q2��r���\���T,<H1��U�pd�+��%��XtAV[�C|�e�۴&eND�~�śC{��"'|����r�B��oF-�G˗n�(&�e��S�Gט��Ù������S��Ef9�E>�}9���vv�P�O4�<��Bo����C�n��K+x��qp9JEt�-�cy��	�C�U<����L�E���Z�s�E���j�I���Y�U4�ˍ����S�EZQ��C7ꌂ� y�D6 �4��,k�D$^o]@�+��IB���,��o�^Xz���[}u�a+��@�g�Km`_����ɝƭ�wJ�+�	E=�)���$��뢊s���p�q���H�* ���}�7�{v��.��i�Aכu�8�L����������ߊL;�6|B����bSW4�w�P?�֚����魖]�zg�x�m��3ӘQf[T�5�AI߷���h�w��9��b4d�n����{��\��z`K��7�cz�ak�^-̪h�\��*z�򏣻劮r�sF#}��}�Ie[�����Y�<�zR�b�������S��x���?��n���܂�l�:�~9z�J.��j��o���JL�V���*|�}%�����xفv�r7^w�����(Ö�=�\�Y��W̧��[ĭ�Դ*p�֋�>�W4X�a��g$�lMJ=�o7�Z��SM߭i9[�r�"Ӟ�]1?�<!�GZ��}O�Cb�S�40x5�ɚbFY%��'���&��Q}�rۃ�R��D���槿et�~(<&��ڥ��6�6�~{��z[��I�m'��c.,����bW��S��(*6n�Q���������dmw.?��[�c!"!�uS��T�K�YZ_�ݘ�O�pF����y�o{	:2�_�"R��i>�\gm:l���8�b}qz15bv~u>�M��|���|��aJ{����1h���vB�9��� �nhয[=���k�p$Dv�2���{��N�-P�2x��f��`���_i��U����גv�l�VM�g=c�h�őP�1�����_y}$��$�%1¶�O�������|o�u��:����lv9W� AuH��h.A�_1]X׻��O4d���*�N/��p�)C���SN�~�����CAt�#�sM��N��p�a����l���>����i�-��S�:��x�|�lu���D��w����~�|-�b��u4�g��0X���n�a�Qr-����C���(�����Hh.N����=�i�>b.�	A�}ĞU�uw�+<[�^���홗�G5'���7O$���W|����I�WS�����J�҄l%�}2ha�4���/W��Ƿ.�.Վ��:�y��`��]~g�Hjb��ԾMRX�o�2�l��ʐ�a���\%k2uy����|��� ���F_���45սO9~���#�eȱ����bj�D�8~h��0��7�a+��xnC�I�������Unu�Չ��m�ʻ���K3�:ݍ q|�/�z�����ˡCv����TZ��ՏӱP�4FZ�;o�WV���҅FQ?��V3��巈�XP�N�y�^//��^u�fus:����F]Z��~"TH�笐A�o�]:p�c[+�S�0	�����p�����;P@�J�G)���.���_��Z�^b��޾�t��a'��m-��]��M@����W�!� �̟�rNcl���L�}'�NrT����9WP{_�����&����������8�Vw�����&�Y��DTE�!$4�[���|l)8�O��<�R�mΓ����(��Xm������S�E�o���ݟ�Z�Wm��~�d�)�[�6��G�%4y���x�6AQn�;��������!`��i�S|���A��gpGVhV�vG�ͭ:s����Aק��;s[���?%�+%ۡV����g��_P�sJy�s$~��M��{T�L����qy��D`P���I'^%��x��Ϗ��<h�Ə��R�]�-*[1a��E:��Q��H��i���j�SJMW/�M�DE �2}�R%���)��֨��4<�(b��4�������)��Xgց��}ZQ��C���~��5?)n���zC����Tg;����9P�Y��׺��ų���ctj-�q�d�}C֖;�n����ݗ���^ͭ5-���8���3I�p��_ۀi�p���#�lw���$�w&��n���~&$O��M��ޛ�j�'�&��dD�{�u��}0�&� �������4HI��T,���&�`�GF<�9��:aK�R���M�B��t;d���c��z�񏥙�v�����;�TΖeN8��e_�Q��}��"�Hn���S#^k˔3��T�ku�dF���:1�/ͥ��&b��כq!j��`z#��k�~,� ��74�R6DDL�%��[�|8��Q��M"zT�k�?S���K"�7ܷoJ��[��3f5F�RJN4�s�7�a�5�)pE����\Pr����O�5��b+��ۏ	��K�9�O�]�Jj6��k*LB�F������'Vʽ�,�5A�{y�j���"�E���h�9S����	�U��9�M@����sU�@ߣ�`*�|�u��!����Ϙ�E"�h���Hw�� �
U�+}� ��L�@���"p�ٔGe�@�^��"�/!�/�on�=բ�������<�,栦��,�Ios�!��x�fFqV!(��q�u�Ջ���Ε(��[I�0�����1����ԗRR)�kS��cu�
��Ȕ�Y=J $O�Z-?_�H3V���]P`N7�1�V�Nu<|��;\�K��v�=C�����y�~>VXs�jʬΡ���}[%����� ���.?hS��ڊ��ۥ�7��3#���	d/ɮn=6z]Ŀ�	�M�A94e%� Α|�ݲ$L��唆��.K���*�V�WoG��:A�ǅȃ�]"�.�ס���R�(3V�z�q��F�;����ؿ�bG�����j�P�\��ڰE�4:�rn@).�L�N�L
���(��'P�)��y*�_Kp7B�g	����L	D9#�7��ƗE�~/��r��p��������>Je��Z�̦\	(ؽ�AR��&x.g,��&�*�ZvM/�������{>�G�H+�����I�� ��I�?kŃ�S�T�����AT����c*����n��}��s/ʜaG�Cn���#\D�(�3���뺘���&� ;�����tt���C��F4��Nەqur�.��ucP~B�wpk$��T��_˒@��"�nP�(�n�:*�3���p\���&H���%�d4����!8��4����N���m�����$TK�~�T�9l`eu���;�f7
}!��.(�X^��i&����~�{�k�QN'�l�3������+J9M����zz�Y.	j��z��On�B�$�Q�� ��B�a�:(���e]p����&��ܷM�ñ�?���H6�t�MFP��Ih��ʪ��Nr�=���|x6)��iȏ��~n�C A5���\�7V0��顦��.8xh~z͑VU�(E�_h7&5�G�P.%NyD�H��6$M"3�t��^p)�2�h];�X3lt����;�R�!���<���3&H� uPOǢ��s=Z���$��拿�Rh���!=�}� 3�(��l0җ
��W��hޟ����U�e,���+�K_kE����q��{����1��+{!.Li��y8t5o=:��Z��y�mo�چ�:"ZgX�?�s�������3�� ���?�Ǳ<K��o��^͊�����%�z�[���گt����/������;�b/���`j��ƒܼ��
ԣ F�������W�G�����8��]
�L{�4�
j�,#K�D	�����9O/*�kjs��/��*�ԁ�c�.rA�&�d�>xc4�����������>��?g♊����A)s�d�{�_$��\^Re`��qE���;�Sl��FD���𫍦��)8�k���ߢ�e��Z0cpnzF��*p�cӐ�Q��x����L�,��_�48���}�2m�7�=�\�7�&$%k�����@��Qm���#���\��q?���ka@�4B�AB"܊�h"�Z�J]E����,��:9M��_2i�x��lbL���h��Gt;�]�|:���Qw��[M9"�4狿��*���җ(D�![�����A ��$���J�LU>ex�׹���t��VK	�(���.5;|h�Q.���L劙�$H-9H�s�<T��帀R��ʬ�}��Dz�n+:�a5xpa��5�L$�� �C��
�W�ϒ(Dg�9�����DG�>�C�ty��_��z��ғnk���Q�rY�@�P��������h @�~� ����Q�g�.�9Qm��v�� ��]�z0I�`��XC'/�7�J��n��L�`S-�)��a3�	����F+}}�YemY� Ue���sR16����|���-^��V�`�|�O�v.��G�sX�<�`�مh}D'���Th x66	�v3��`H�)���8���K
����!�h��	ZNHYsC/��m��/�Xﰸ7���b6ɝm�4��x��\J��-<S���v*��������X��~-��.��%��D�Y��<X�$O���"�mT�b��#꽟Ӂ*�;�p�@u�K���B��[���]ˢ�.���[r�����o,�J�`ْ0Y�:gg#Z�_�3t�{9`I���^��������?Y<9�x>����1���
�92��H׷84��}�?.�J�(�������xp�q��76i_�H�ʽ������S3h��[L� �j�WG����õ�=U�u���h�{G��Ԋ�u	ae�/���;d��X����9|���Y�� ��U��q�/�2F�(��Xm��N7��-�Wy�{����tr��g�kb,�֚Ƶiz� Q����`@�{\�U���wx�גM%���v>I�d�/=����Ջ�oy	�o�5��٢����*�QT�G3Zw���'����7�2U}�qu�����smD6��cK���G�$�J0�VQ-����Ƴ1���6�\_���M��b.#�[�����'��$$,������>Ė A���ɇ&^RJ>�L�����Ȭ���g�+d��� ���ʌ.5�CX/-�1��N���5K�i9�4"b��V�ֵ���!�QL�����%�^����(���>�=^f��x2]�#���I���
��=��Jqf&�j�4K���m�U'� P�ؗե"$͓���?Ʉ -0<�-KY�M$��56H����������p �?���Wb��ݻ��+�м^;N�j|��H��x���X&�	:��"}�%_E�>��n�?j��8��&��H)[ �i�M���~e���E�4�Qd&��
<�Pw�Q��عV����(�C�$���XT����Js�e�ד��j�vx��B�[�LZh�^�T�����dyv Jx���OW��'��*��^6�K26l����|�{Odn��6�zs�Q tT��x8�J��nӐp��&:���9��n�&?.�:��p���� d<��J8TPR���.)�r�zFyO���@����[Q��*�'�T!Lڞn���ཿ�egQ��J�^Rz�;�~ĕ"q�_�o���Y�`5L>���`�S��^	���t�?27�LqGJ��������2j��DJ�G� !�I����˓�I��f��wn��倾>Ijo���M�
0ğ�Ʈ,��Z�4�XٳhmJ�V��7��Z�>A���	J"j�%���:S�,�@���'�۰�> �H]�e���n�Zf�"���৊
L˔�d��/��k���Z?Eo&2��L>wr>h� �8~36�dt���P1tXF(��I�3�C�K�ۥ�{�O���>q=z���Ķ_�M����ޢ������9��徊RިP�.B�^�ȩ�l-Yȼ��@��(Ǿv�LYy�F.�1d܈�⧀F���M�H�m.���ӈ�yu*�be a�	���H��iȀ�a�s�@��?�6ӳ�MP!w�8率�gc@%�2�g���*����8��i:]�r^��]�%FlB��ms��֘?�nu�y����V�'��� ���wz^p*;Pa��X�h(;!�Sh7[Yc����Y�H���P~	�ΎK|��L�_[Y?&ᯰ�"⩋RPZ�}��<[T��J(|�(څ	
�K~��!%��%В�=`27�IB|��)o� �:"@Ȃw����������j�V�õ�����膶@�*�/Ĭ�b�<�AU&���o�](W�T@!q�$ܯ�2An�S����7��ʴ*��T�Zf�����}�J��wu��Į2��M,��t��HJ:ǃ�]�yj�?��E��~FK��=6X�	�YD]����1c&�n�oS���Z����Sޯ���XԵ̆Y��2�C��Wq�߂}kI�U(d�a7�q��I��>oj�����Ta��z݀�-�D^��&Q�<��<�.�A�q�*_��	�S��$���h'�GP�$�4��������c��}�A6=F�[cL/,��_S��=K@n�+.���W�px�qt?�W_Z2����_�Pv-Jz'c$��0U&�!�'�\Y����a� (��Ν�A��1*���v��l/윎Z��?�A
���e.C�z�x�Ԅ��c����;Qs@u�77$�RR�t��U
�
>թUY�W�����_��O�nP��]�xT__r�~P��&� ��ݡ�o';�����( ��k�DiB(�I��0�#�K���q]�IF����������f'�#@⺷�j��ɤ�/�F/aD��q�v+cZ0�{��m��O�Hz�JVy)ԃ���D���(�����YkJ�,1(�!\�Y��ϓw�8��ä?:\J��"UQ.B����c|E��/��qj�X7t+��%��W�9�U�������iZ����{0!��ͧ�c�� ���M�P��ZA?�)Hfm^���ya7�"�(���W7K�}���♐��%�
��~�<j����2+u��Jө�kq���/d�/h�D��7\D��0�6�
���Tn|x��#�ݬ�0���T��#�	#��)P��ѺC�;��TE`��,@���X��v��xcu��Z4��;���=�]���iv�	�k
f^��{r�>�J�ܦ�w����4qX�o�q�y$�adF��d2F8Z����k��֝��l.GحLm�����$��G|��������l�e�`�Q��Hi<d��5A�U253�]QAB�z���A��2>	q �3nq���ϣ^��C�6@�ޓ$!�J�f�{��/}p�uֲpN!���C(��B)8Z�j�!�"|�P��-�7#$����#y%�zwZ-n<@�j���<7�>͛v��k�������a�}�q���췬�eA&�*R�BȀ���hx#tWI�DmS/�̄��M�R�`O��zx�U&���I�ފ�'H�bu�'"�|��YA@6M���Uix��2�� � xv�/hN8�o@���di��
��k�Φ����PW�,�^Tn��B�|(�}��3օfm{|�T���~���!ܸ\����W)�(X�{<4\�f7�+�d7VA�`&0#�����7B���J�LbO��;�{H}- ,ۏ@�d����2��v{�	s��d�[���j ��2����R�C���D��$!�~p
ղ<������j�x�� �fl4��4Y�E�b�A�*��%P�/ޞ��,��(�����B}:�[�F��/��HOp!�G/���t�n_����!,�����E�/��8���[y��VdN|����P�p(��ԋ�CQ��}����dD�3�?&�e,L�2�:�9�?�9Nؗ]o�|}���c�(�1��o���(r���^�R�a>�=^�B\���$����@�����r�\��<�畉� W/�y�Ro��0O��0�Se+BR�o�P�G	+UL��8�H�K�;�'��'k�=^뵫[Մ��(U�&�F���@��{:��d$�8�qI4%-�ԌhwP��f2�b�956�?�h:��!�2�@W�Mu@?#��L�b��_V�И��Z�ia��q�ڇפ�Q6+���[}��	#4E��B�(�j�m���<c��mOߵJ��=���9m�C
e���7��h�q"�$w���X�P�e?W�(���kY�O.D���~BVܵ���O�L7tq��s=�'�xCTz�/����
�?�WR5���A
s���������OU^����I��R��_�_���f݇1s���Z	{[رbK�D�����Ǳ���()��40������+�፲���N?��v#Y��FSVA�`+���|?k�9[�%��:��H��h�c��и���;X���*��9�?V �^�]";�n���0�bx��'��}e�[���:�UI�-��$���}\��t�� ;�k?/x�{!f;�C|��)�¤Djj�݁���#W���/�`Π�Pb^5>������!�]br���VfC�"�c�O���fG͹i���7kY1�r ����A���(�h�K�qҧ��N%��ۗ%Q�x�)к|�ڛ�*Hg���N��3��m����PK��"R(�n&���48��\}�2�W�Z�jW�� ��������&@s������\p�����'D͉r��2�)�<�-�f��]����x�ĕ��pȸ���i5]Hr���e�M��%��EoTkL�������PPhv��Xy!�Vc�ة���'�-�a�"y�zp�R�M�f���̬I���[i�+ߩ�Yf,�71����K�5�>`�����|����P�*�����_rXȡ &"oAL󳖂60⤭�֬J�@:����ޅ:�w���`�|:�[�~e�E�P�_�s�����c�0���;�3˽��N���[�����xY/ ��C���.��;D2�ܗ����8)�-��+��B������V	-��C�V�G>��2���6����Q���2Q~ۇ��Z��z��Io_��pl��.�b�VC,J�%���Iqf��+�򒙓��1k�ζro��0�l�bD��ޟ�g��&��+	ƹy�oG�������]s��PMT,��p\��to6K ~�?�����Z�u�N�H�O��&�l%����:�3>�������ʬ��������I��*����R���tI�^����Q_��~�$K�$>����|���������"?���6M�ĭ�GD���Vtm
��V�6#�B�No�N���;I�@{"��J�%O/�j�cnF;T.�q�e�E0��i�@u�k@�{�
��o,2���θF�f��s4eD�'�&��"`J>6�Bb	QOn�,>�NR7h@k�h�A�d��������QVAbe�i\��c �*� g����:H�L��ۙ�d;'�6S�C��px���E���|��V�$�GE$���A�2va4 ��1-����@� ���(�Ҫ�7z�䠁!�(@����>jK�c����H��ȝ�~L�:,f��s��>��� fV5ܭ����X��@���¾#~�qH�g�z����X�pй�r�������� xIN��).���ݡWst]� '��LZ�p��e� |���%^G�>]P��!���t�;��q2�|��(�ɍa���0S;."�y�k��*�c�婁[��c��t��H~���������M���{T&M�K�)��y�&���Sd��|$���{�1���c��/-�S�t��/N����laU�//�����O�;� z�)8{(�n$ͦ$��5�P+�#Z�k�����׉�ѻ�gm��j��ʷYs<��x��ϳ\�Ý����q=��jF�l�߈��_cSl�Ai��c�Hm�t�U��~��:��M4|����o����ř�r��H�f�_�NY�HZ��^�H�Į����ĭ�f���&@>�5�z:hR6G&�%
��
���LY�[� ��V$g�U����&!b��[�X
z.#,LVu�VQt��u؉k (���[oiw�}[������鲞����@z@��'w*.*�ԟ!�x*�hdoct����p�(-��nb�*�)�ko�O�v�o� �#�3�cv������j�'`v�cz�N�=״A��+�ol�C�'�N¦��9��d�����p
N(�&�����ɔ�@}�l�t��j��n/MZ�����-�D�=��A�;^�8�W�^�U�S6k�j�p�V3�>#�ldC1gc�.�p
N�-d��
@�a�v�z������c����fQt��N����E-�i�K�;�>��(J}�R����2UL*D,�C�o���o��K8l�-e06/�A���8q(�]�4G�!��VN����t�
����H g��}��8j���P�tg����(�i�p8�	�{k��2D%��2��%��q||�s��Ǫ��iXK-k!NƆ̒Y����q�"xUP��M�Q,�^�kϛ1u� �д)�,�r��	6�FQ����$q*� ��_� 1���)�?��uD�X�?;˔�(�p���XG�Ƿ�=���L�,���APP��g���_!t�=h7��9oP-��z��3����޾���C{E0=���̆-���?C�6�N��V�,�8g�.#�o�>8��SGCo��k2:Qo�ͳ��/.����[zX�G��A	���x.�K����΄���Q�X+���{#��@&p���τXVAko���]b亍��d�%8���,�������U"r��1CI����(B��%�<~i�؀"���>�Xd $�R�Z3t\l��&�s�־�_�K�Z��rg�[�#T�ex����a4�a���9	�2�$��ʠo������}�4<-��"�x����G���mi|g+�3F{���C����B�*Kp%`����>q��2�P��Z݅�ޚ��0Pր���zD�_X�_�S!�ޮ�.F1 "��ᢶ���#�nɿ�.}�H��R�=�P8f�) ��,���}����u����?��V�̎���Nm�n�9��[	�� 珆�Nu��.>��Ax�ϵ�g�����:<��I�Ezj�Q�{�N=���o����A�o?�x���i�-�Ȼ��]&˶7QE��e����s�����=b�I��Ό]%�j5��l�zL�����p�.cv�̫R��jُ��,��"hT����a(���R�C��1WZ�~�Q��	őFt<����|ԇ�(��X4�g� w��	+-Gq1r1c�Y	�,�*��>�a�̰P��(�ۻ���=�PtR���1�i���&�g�G��$�PJ6�Sg|�:���,�|�CC>���iM	)Z���Ƈ�W��h����j���Jc�xk��}�8�׼�T�G)F���P���b�X>�g���)����5۝pa�������(��Y�'$
!T��"���B�mΟޯ|�i�Ò��~��L��8���PX�z�\��Ì;�=O�4�;͓��:����#�#��Fe���M��r+�o��ʹ�*0׫���"�#}@zm���k@����:&�֟-xGC>��y݌}�6��5�w�c�^|��S'�kA��<�9�1C+�.���'�W-���,���Ycq�[���V�S����j���G72m܆�NqÜ}�8*i��g��t���#�o6�$��ߥ�ҿ�v|'����J)%��ul\nٛ���ei��I��Ό���n��G˗:�Ai�#�f������}*��!-��w����ާv_i��q���v����GG5�5�>mΞ��K�?7��{#N"����<��E^.���;&��<�-ԌVvl�PM��&��S�����˨~��d0������֕`4*3�2F��ʤ�mv�aN��
�#9��7����*��X�F�M¯@C�&�iA'��j̝�s��^�|�{�CvC�=|s��+|�]�;_>_O&J�Z>�5�&�F���nH�2��p}<�|1��{��&����|I��3H�!��y�|�cM�l��JlYl�D�3ϔ��ji������;;h(��W+1��� PK   :Y�h�F  A  /   images/cb0ca54b-1964-4771-904a-f612fb73280a.pngA��PNG

   IHDR   d   �   �8�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l\�y�]ޗ(:���D�uR�]���ZM]'q�&��Z>MѸ��nݢ���h�(5Ңhc;��I��)Ԋ�;�uZ�e�A�(RI��!^����f�����ݷ�%�����������̛�.R�N�>-����|"���F�'?�Q�Q�P�J e������Y����Ν+R�R���f ���CY�R#l 
��栣(�d�䠔�T��P�Q���쓨���S�NY�
0�b�"	D�(KP
��Ԁ,�.U:A"e��6�W����;�υ-M)̄��!���r�R�La��!n�u)�E��G�e�Nu��f� a��~�e/�m�GY+l�C)���|$a��g:�WP.Cy�޾� %��R!�X��Ua��!�D"���;7==�ppp�J�7(lp��	�P2�D�e��m΄��T@����j�?����v��/;;�6++k1��j�p�B�9�4`(-��+�mg^Gi�'�����!��7����P�B~ p@\�����<���,����������v	
�`�8((��By���K&(I�F�ߊ�u"�TXz_cTLDЇ���QW��S�%	sQfARN���!hi�R��w���k��`�@I
 
�RF]X0�0������򾾾�J��q_`2|RQ$��?�/��f���~U֪���ɛ[�5�y}2@I8 #N�&, �,//o%�+HKK�����TH[˽������C�Q�B�9Ch%�{�\	`�AZ5o�@�o����q�Ii�3g�H%��-0���*a�'dLL�����9�R������Fn�D��^�BZ �\x^KQ�0*&��b���dwww柳A�K~�(]��sJ MMM֧�\�ޔ3�d�nڴi+�>��E7� @��P_'� ŧ�E=' -�_�e��KbІj�' �>))B�üٟ����`"UW� ��+�Y~��(���������`D�$(��:�٦4ؔ�s��m�}/��"W���H�$��36���?J�=I l,T��{ɟ�
۷�� �Tfff(0FOS2��� �-������`��@I������7@cIj� �t�*�&ı6� J��H0hDi;�D�Ҁ�a�&.��p�z)xu�ۼhA(Ð�Ϡ����. ލ���죇��!d;i{֡��!%����R:�
����-�)q�pF"��vآ#^������ǌ{4)u�t��e��H %�ˢ�\&�G�A��Z����d1j��h=F�P�6$�=T�hX7U�<L�ざ�1{�l��9 Z�ragnu��4z{�A��{dl�O ���!0N��H����M�)����r�v�3~b:U'	Ƒ+QJ�12��O+�-h��)����(3`?JEd0Ҡ��(��~N+�om�� ���<�8Q6��8U @ F��v&�N�� �����2zO L5pzTg:=�l&�Dd�*�h:Q�kb���j��-�N�d���TW ���l���po�&$v��}�3VC���-���c�AxV�rb*l ���f�#Km�Or���5�y�#��v0<��U�*�m�N�'��R�"1v��d2�G?�y'@�$�ľ��ūJ=R �X��Q�S* F��:�`؏sb����)�W���� ֗�<@RB�����>19�6Dx��z�������Q�j�'«,b2$�?�@��׀�"��P��'!y:�&|��F�Q:<�T��K��]$�� ������G�\��2�Fi��dP� ���Pτ�I�0hJCo�R!c���2MC�c�	0��w��ܹs�>,���˗�[TTt.�{�K�\%(<����͚։#���b_III�b`$"��������Pw�yԓQZZz�2u�����9s�����&��E~[ОN/���HT���YgϞ�&^�:.���z����7�p�OM����*������;�g�dnNN�������q=��f���C����RH�d҄ �tww��LɄqB��>|����� 62�t�۷�#T=`��]�v#%���Ou���Tv����ӄ ����ϥB!AЉ�<r�Ⱥ���c�����-�8q��<��+�k�׬Y�*�U'�R��n����h׮]롮���l����
�����疘#����������X���P\��+�JJ�����U�V�����UIA���ر�؋҉�j�Dܔ�X:P\�ۡ� ���~
	;�����ח�}��o��MJ�E�eECтH0�����ת���@%Y`Hg"c�֭�Am.H0H�
�h� .^���%K��\�f�AW`|jsq*�A�Ҁ,Z���+V�V`(7v˖-�ttt,K50HS�*؋M�W�ޮl��� _�W�:� M9@���!z{{���!�AzT۶m�bkk땩�M��)��ٳg7!
�@Կ����:����������SҔ�`̘1�F�A�5�cj����G��"�Ju0HS�Q\\�VSSc��"y،�S�N1%R����DQJ��,gB���pm�+Um0�R������X��p�ڦ���@B��6����333&�|0�Cpoi��p�|s�������n���P8<<�'/��&ـX�|�dF8�O�����j2�!G�O�!���!D���`P�>���Ո܋�j�>�*���#ZJ �_ �����`^V�s�PF���Ա�)Xǳ�֡���jD�"77���3sp��(�|�]|����J �� �<t�P�{Lb�kڞ����pFv������⥗^��w_\7L8 T��W�S'O��?,��]UVWPP��i|
������r���'%e�ƍ�{��~	�#�r.>�`�'bB2���6m�g���*�3�������ӧ��1�Dn>�\5tp���'�����Z���~��и	� 1@^~�eq���t�D��2�����{'9�F`K!��)�� w�À�}��v'�$�2��@��#\NI�/�[}�E��^��B}����*%�B00�
蝰�SD2tb�Ҡ�+`۵�x�߻)%��b��S@�;�(�{�d�[�6�n|	ݘǿA\����?��},{
Hvvv�5�z��!�6�a�9�"ˠ��u��W^yE�u�]QU�) EEE�����%�ħ��A<���ܗ����3�׃�ak���s�Ԉ��x*��Ə{���ȵ`QW� t� ~�c�S��;�ݬ@��]�������`!~�ɍ�s�C�Z�	�IM!�m&m�9�D)mg��A}=Ѷ�3@�2`v6DFtqqsNN��`U��r{
k�������p�

��nK-��]j�	ڕ�X���J���y�e��8��n�v�W[[{�}�ܠƗ̇dT�*++���'r��\�s��JrqG�X�Z�r��>6௮�N�w�[9;��?�ݗ7�f�D�ZE�w�	rcL� Q��3@`�Ekk+|Y�F��������=��Q�� �8��uww�#��]W�)�t�j�c_���,..�_Q��i �iН=S=R' `8gA������?%rY�R���(AHI�ta��k	���� ��%��\�pNC�ma������%j�J���7�|^2�F�1~�����|	'n�b�����KP T���+w��2��+�3އ��+��#��P�����w���:�NL1W���t��"�|�^6-:{�,Wd�1����ӧ��+`�4�Ch�BF����"� ��\���G!L����l�(ޅx�G�2כ/���p�677gp�u��f̰.e��,U"&���Ioii)I䫁"6 N�"ҲS�:�u���!��h�P� �/;��C!Eڒ�dS�����`�w���b9mkW�Ĺs�Z�W(G e�	��C�����)���-�����xYYY�+k�
�O��h)!��!\iB}ʆ���q��:TU�(� D�AG�����FK��p���%%%�)��ȕ�#_�4٤E�?��������[�pa@�G�l'��9�[�lY������Z>Jܳg��3v���+�.�:T_g���5��KOO�80�@���a����#q���6�F|޼y|gT�����������j1s�L���'�M���lc	��ɷ`/^��H0(8�'���ӽ�1��V��Q}=zTvl���V�8��QGP��SlE#7}���TQN��g$���P��s8��P�Z�*�x���a#KKK�r�������5���JUV�	w���yZ���}qD0��MqX,� 8�k��>-X� ���L
���!�>�G���*P���:�w�^��c�´4�����܉Ɵ;�Lc�M�^$iN>h�l�'��?�s�Μ9�O	vzRtH��<z��!!�7y؉�_��+W���M� d�Nv���.�@ 0���lV^^nƎC�1�Q��j�Imܔ��+U敽����ol`.j&�s9O&�����Q��ީ�N��`(�
;$r��X�U,+Mt�fԎ�,��!JԙF! �+����DG谟#T�s�q� &	-���rb:SU&Y��z��ĲzH���}0H8o_Ku鳉�ca�y_�LZ��S/�r<4J 8��B�z^K�/_�N.Rd���_�7J�dHMM�%��N�q����������3��t)/��u��VF�M#* �-}�b#U�M���7N3U��
tvv�.�	DEE���@�X?�Ƴ���J��X�"nz��-�Do���>����2��%K�9�#2@�ljjb�����f�� (d�Rj�˵�K���)|ǭj��)=A+x�4�  ����H�=0A�A��p��=���</O�� 
�N��ןm\�f�ZF�A���F���1J9���||�ɓ'-L���[ޙ
,y��A}���.MT{�^�S�Jq�:�������WI`�g��|�P����ӳf�=N��<UY���v��|���:�`0A{sJ2��5�L�����Ĭ MT)1��g��ըU.�ܓק�7���) �3�K�:7�z������	��G��=��hԾ���Y�ٹݻw[^�ڵk-�n�)���8.�P�%�HWF^3�]�0��|T��|��S3}&�;�cǎ���F���4~za3���>-&p�֦M�,�N�F3R�G�D�p$:S.\�$B�,�$1T���ie(��4�6�^RR6�$#�:c"��@���S�Ȯ��OR���؉��� ��&�9��;Y��$s'KZhP?��+��t��~Ω�ɶp:ٓ'D�A�8g`�D	%C��Mi<Dُp��a$�m۶�֭�s߾}�p�6�������^��5�F7ʧ(o"p�T�|�����G��m���i��$S`l�^|�E2�=0`�jx3w�Ӻ��.���� _�}���O� PJQ�;0ο��ߢ�?���/\��o�P"1�?w�Xr+
nIэ�C��YpO�g I7U�CxLzL#`ހ��Dk�K��x�[wL��h~���;<�͌x����~�j�G}��<DSW���Z�K���ׯ_?�]|W��H�6��IJ�Șb�7�x�/�S���xb�������:R-V�5��U��|��	���mo�t
�^�-� ٰa��N��K��hW���BOS��!�C۷o?B �9d�Ν;9s���Uu���=d�n�&�������x	J"�M��;�K��mLCu&�� 	TS,,�z5�@���ǤeY��~�l��*��Q�N��!y�ózF�/�w�M�qUA����#�Wop=�Q�\%��_�\_.��x%%q� �N��4���0�P���;���3A����(;Be�^[C0�m�_�?��m�ߠ���/(q� �P�����E��k�?!K���wI�ek��;��Ư��P���xA��(?G���h�)�#D�M^;�;aK@8��Sn��^��h�b��ⶐ�}~]�eyh� 0h�~)�����fV�����r�N�1<�.�\�R�r6w�i(O܋}'�(l� fP��ghh k/����#D�9���a/2���0�i��Ly���ۤ��i�?AYcp?��-y���g,�DH0�)�F�\ AC���_6�����BuVch�<w�K}_ $�r��l�G�L��d�1�b�����u�Z�b��?l}j%=�?2��Ca�7��B5�D��3�<#�x�	������-۾Q������Ai�h@1���h$���(/�z㴀�{LUԵ)����o��C�O&n��;T׏���=!q�*PN�)(�����h�����G�F��+&��������"�)u����6�A(�(l�}�0#��nQHJD@`� �%����^�e�\�hP�dP�~�ԱGyD��M^�5�z9�Y���t�ե=)5l+��"�nR�v%, 0Jeū�9qt�.��Q|��p�`^�dA�"z�5n���m��d�c�=���S�t�ɋ/�������JH@`p%;e��)bҐL�V\D�&�>���{"zzW^�KJ�m��O���~�m��m ��CJ�5��qLp�ѹ��Ы�9�+�N��������3�֧3�v��%l�����Yؠ�j��uy��e�8@40�8�]�����
��-�@8�i��f��/E��k� Y#�r,��u�B���S�J^�"lUr��@��(�
s�'l�oV}oξ幜C��k;m�-���ʗm9�"(xTC������p�?
���P��8�7ܐn28�j0lt���%�C�Y���g��5 t��8�}�����C%]Ј��aN
�&���D�0�O����I5L)q�j�&׭�< �<�A�c�a~�Eqq��5u٨��:©�
��l�A�'�s*�ݦ&A\PhS6�)hI��=�4��\�C:(B�����%]mp��L�H\�'w�`��r�۴ô~(T����A�2��m!Ϲ(ĪG��o{%�	�ø�ް�2�;�{<��C�a�8Ki�s���
�쯢�/�Vސ�	���Q@o|���̴���]���@̰����wĺnw9�m����T� �s�\˕w9����{�+@����$SѣL�c��3�&����ã�ئ�B�~Sr��W��,܉�g��$]^hB?�!m@��쳣��"a��h��z/E��^�Ʒ,�鹲mGb��s�B�F�;�r��G�za��3��7����i����^.D�u���Ƕ��M����C	���z�D�ɓ�t�E���U,08�db��:ݖUxx?&69��s�����ɢhfo_S?�QZ���9&�'�:M��RB��̹��% ��Cu#��d3�3�{2�ӓ�"5P8
�C7@�'�?�S��)��{�H��s&�N2i[�d�t�@�%1wo�mx����ݲ�R�P���|�I5ZM���lw5MJ��=���~�U'��v_"#2�c�_p�\� )F�H"�~3�$���u���v    IEND�B`�PK   %:Y�2v�E  �&     jsons/user_defined.json��n�8�_�0�;��N�wJ��4�8iP�
J�al�Ւ (�@�2�LCYv�X�B�̍s[�Ρ��\���a���aU��[��$��p4��y�d�� �p�̙�
�[�������Z��~:�N�*�'��֩.�<Y�����y�c
F`%Uh�)�".@LDZ�H+8^�7�$2�������x��
0�U�f�J}��&��YU.�rx=ZU7]7�ռУ�2I��8N~�o���4�^������4@�y���<+����dnN#6���6��.�F�{ �ИAq]N��m�׍5)���2W���u40�f������㔐CF��٤f�E�Tڕ~9'���M�u�jC���".I��I�Jos2�.�ӤX����l^Ԣc����4���Kt�0Z]2}�Ar�ݩ`^�7\��R�e��o�l�Tj�˚�;e1G~����N!���i�r��mv�����:jF��"�Cn���{��54u?��Z�U�²�u�4���a��ܖ��7o�4	���0��b4 ��P!� U �ǁ XB��Ӆ�Y���j�j�(-ԍ�����y;����Q�-n���(�|�aUa��^[��Ɖ� P� H� �)4"1�"�!S���8Q���р�$'�����8\��� ��c�:(��p[���\PocsJ��Lvp5���1}P��(���|4�G���ҁM�&��{���ݞ�z2�f*�1��#Q�y���$e��6�e6���C��d��W'm�x�:e��eu�z���!|Ww�ȵ�D;��j�|pUۜ�ӄ舍�S�g� I�i/� jf!2�HeB��zR�a�{G�;��p?��$��f���
�������\��$���֞�d 	@TD003Dʡ�_P�zL��^`�`,���f�D�f�j�0Qw�$m�x�-*�#Um6�X`���v������"����L���N�`� ;�0�3{��:F�]]v�cl�c���S�>��Ǯm���C���<���*/��:��K��tU�VuϮ.\Յ�x����K�|���zv�n]���&��wP�
������c{�t��E�������0wp�0Wǧ�m�y��8�Ƙ��M�6̼�Q�+{�6ϼ�S�v�q�h�߫}�!�6Ӽ�[�v?�m�yo���nS�{;�o�ph�۳}�X��XvEٷ/�pɮ �vW�]�b�ώ>�#tQ�
1�����(v7mrp�����M2݂&�|����y~�;��<���J��V�jҿ�WGk҆�/敵Bpܿ�����'O����j�e�wr�Z�����*`]����z�����ZP&S�*i���p� ��'���Dz�������c��1�>f��J����œ���:,smN$�)�����r�ĉ����ö_]��$��R�@EZA
�M=��ʌ�����v���0f!�R��8�fDT�,B4(Z�M�f&3-��[�znfR�.s1��%l{�}U}w>�˷'Z���G�c�ߞb���g�/�?ۧ>��U� ���-g&�#��eZ���8���]��Ex1�yĀ���x�o�.e�t�9�~ِ��PK
   %:Y��+%  �g                  cirkitFile.jsonPK
   �a7YmS�;F� � /             X%  images/45855a06-4846-4a51-b2b1-60b9838f281e.pngPK
   �a7YN�v4	� m� /             �� images/4949577a-1080-4c93-a0f7-9bc81c12f32a.pngPK
   :Y�'���U  �U  /             A� images/79f1f6d5-8698-44f6-90ff-b688d5ed2669.pngPK
   :Yd��  �   /             X� images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   :Y�]��N � /             n� images/907530ff-a8af-4c9a-ad67-f4101e76dea0.pngPK
   :Y	��#u } /             �K images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   :Yԯ�|�] n� /             � images/a794cf5c-4b1a-47ff-be53-d48f5d14bb41.pngPK
   :Y�h�F  A  /              images/cb0ca54b-1964-4771-904a-f612fb73280a.pngPK
   %:Y�2v�E  �&               �= jsons/user_defined.jsonPK    
 
 j  D   